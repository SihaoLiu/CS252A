module GPA1(
  input   io_x,
  input   io_y,
  output  io_g,
  output  io_p,
  output  io_a
);
  wire  g; // @[GPA1.scala 17:16]
  wire  p; // @[GPA1.scala 18:16]
  assign g = io_x & io_y; // @[GPA1.scala 17:16]
  assign p = io_x ^ io_y; // @[GPA1.scala 18:16]
  assign io_g = io_x & io_y; // @[GPA1.scala 20:8]
  assign io_p = io_x ^ io_y; // @[GPA1.scala 21:8]
  assign io_a = g | p; // @[GPA1.scala 22:8]
endmodule
module CLG(
  input  [63:0] io_g,
  input  [63:0] io_a,
  input         io_cin,
  output [63:0] io_c,
  output        io_G,
  output        io_A
);
  wire  _T; // @[CLG.scala 18:18]
  wire  _T_1; // @[CLG.scala 19:18]
  wire  _T_2; // @[CLG.scala 18:18]
  wire  _T_3; // @[CLG.scala 19:18]
  wire  _T_6; // @[CLG.scala 26:21]
  wire  _T_7; // @[CLG.scala 26:11]
  wire  _T_8; // @[CLG.scala 26:31]
  wire  _T_9; // @[CLG.scala 18:18]
  wire  _T_10; // @[CLG.scala 19:18]
  wire  _T_18; // @[CLG.scala 26:21]
  wire  _T_19; // @[CLG.scala 26:11]
  wire  _T_20; // @[CLG.scala 26:31]
  wire  _T_21; // @[CLG.scala 18:18]
  wire  _T_22; // @[CLG.scala 19:18]
  wire  _T_35; // @[CLG.scala 26:21]
  wire  _T_36; // @[CLG.scala 26:11]
  wire  _T_37; // @[CLG.scala 26:31]
  wire  _T_38; // @[CLG.scala 18:18]
  wire  _T_39; // @[CLG.scala 19:18]
  wire  _T_57; // @[CLG.scala 26:21]
  wire  _T_58; // @[CLG.scala 26:11]
  wire  _T_59; // @[CLG.scala 26:31]
  wire  _T_60; // @[CLG.scala 18:18]
  wire  _T_61; // @[CLG.scala 19:18]
  wire  _T_84; // @[CLG.scala 26:21]
  wire  _T_85; // @[CLG.scala 26:11]
  wire  _T_86; // @[CLG.scala 26:31]
  wire  _T_87; // @[CLG.scala 18:18]
  wire  _T_88; // @[CLG.scala 19:18]
  wire  _T_116; // @[CLG.scala 26:21]
  wire  _T_117; // @[CLG.scala 26:11]
  wire  _T_118; // @[CLG.scala 26:31]
  wire  _T_119; // @[CLG.scala 18:18]
  wire  _T_120; // @[CLG.scala 19:18]
  wire  _T_153; // @[CLG.scala 26:21]
  wire  _T_154; // @[CLG.scala 26:11]
  wire  _T_155; // @[CLG.scala 26:31]
  wire  _T_156; // @[CLG.scala 18:18]
  wire  _T_157; // @[CLG.scala 19:18]
  wire  _T_195; // @[CLG.scala 26:21]
  wire  _T_196; // @[CLG.scala 26:11]
  wire  _T_197; // @[CLG.scala 26:31]
  wire  _T_198; // @[CLG.scala 18:18]
  wire  _T_199; // @[CLG.scala 19:18]
  wire  _T_242; // @[CLG.scala 26:21]
  wire  _T_243; // @[CLG.scala 26:11]
  wire  _T_244; // @[CLG.scala 26:31]
  wire  _T_245; // @[CLG.scala 18:18]
  wire  _T_246; // @[CLG.scala 19:18]
  wire  _T_294; // @[CLG.scala 26:21]
  wire  _T_295; // @[CLG.scala 26:11]
  wire  _T_296; // @[CLG.scala 26:31]
  wire  _T_297; // @[CLG.scala 18:18]
  wire  _T_298; // @[CLG.scala 19:18]
  wire  _T_351; // @[CLG.scala 26:21]
  wire  _T_352; // @[CLG.scala 26:11]
  wire  _T_353; // @[CLG.scala 26:31]
  wire  _T_354; // @[CLG.scala 18:18]
  wire  _T_355; // @[CLG.scala 19:18]
  wire  _T_413; // @[CLG.scala 26:21]
  wire  _T_414; // @[CLG.scala 26:11]
  wire  _T_415; // @[CLG.scala 26:31]
  wire  _T_416; // @[CLG.scala 18:18]
  wire  _T_417; // @[CLG.scala 19:18]
  wire  _T_480; // @[CLG.scala 26:21]
  wire  _T_481; // @[CLG.scala 26:11]
  wire  _T_482; // @[CLG.scala 26:31]
  wire  _T_483; // @[CLG.scala 18:18]
  wire  _T_484; // @[CLG.scala 19:18]
  wire  _T_552; // @[CLG.scala 26:21]
  wire  _T_553; // @[CLG.scala 26:11]
  wire  _T_554; // @[CLG.scala 26:31]
  wire  _T_555; // @[CLG.scala 18:18]
  wire  _T_556; // @[CLG.scala 19:18]
  wire  _T_629; // @[CLG.scala 26:21]
  wire  _T_630; // @[CLG.scala 26:11]
  wire  _T_631; // @[CLG.scala 26:31]
  wire  _T_632; // @[CLG.scala 18:18]
  wire  _T_633; // @[CLG.scala 19:18]
  wire  _T_711; // @[CLG.scala 26:21]
  wire  _T_712; // @[CLG.scala 26:11]
  wire  _T_713; // @[CLG.scala 26:31]
  wire  _T_714; // @[CLG.scala 18:18]
  wire  _T_715; // @[CLG.scala 19:18]
  wire  _T_798; // @[CLG.scala 26:21]
  wire  _T_799; // @[CLG.scala 26:11]
  wire  _T_800; // @[CLG.scala 26:31]
  wire  _T_801; // @[CLG.scala 18:18]
  wire  _T_802; // @[CLG.scala 19:18]
  wire  _T_890; // @[CLG.scala 26:21]
  wire  _T_891; // @[CLG.scala 26:11]
  wire  _T_892; // @[CLG.scala 26:31]
  wire  _T_893; // @[CLG.scala 18:18]
  wire  _T_894; // @[CLG.scala 19:18]
  wire  _T_987; // @[CLG.scala 26:21]
  wire  _T_988; // @[CLG.scala 26:11]
  wire  _T_989; // @[CLG.scala 26:31]
  wire  _T_990; // @[CLG.scala 18:18]
  wire  _T_991; // @[CLG.scala 19:18]
  wire  _T_1089; // @[CLG.scala 26:21]
  wire  _T_1090; // @[CLG.scala 26:11]
  wire  _T_1091; // @[CLG.scala 26:31]
  wire  _T_1092; // @[CLG.scala 18:18]
  wire  _T_1093; // @[CLG.scala 19:18]
  wire  _T_1196; // @[CLG.scala 26:21]
  wire  _T_1197; // @[CLG.scala 26:11]
  wire  _T_1198; // @[CLG.scala 26:31]
  wire  _T_1199; // @[CLG.scala 18:18]
  wire  _T_1200; // @[CLG.scala 19:18]
  wire  _T_1308; // @[CLG.scala 26:21]
  wire  _T_1309; // @[CLG.scala 26:11]
  wire  _T_1310; // @[CLG.scala 26:31]
  wire  _T_1311; // @[CLG.scala 18:18]
  wire  _T_1312; // @[CLG.scala 19:18]
  wire  _T_1425; // @[CLG.scala 26:21]
  wire  _T_1426; // @[CLG.scala 26:11]
  wire  _T_1427; // @[CLG.scala 26:31]
  wire  _T_1428; // @[CLG.scala 18:18]
  wire  _T_1429; // @[CLG.scala 19:18]
  wire  _T_1547; // @[CLG.scala 26:21]
  wire  _T_1548; // @[CLG.scala 26:11]
  wire  _T_1549; // @[CLG.scala 26:31]
  wire  _T_1550; // @[CLG.scala 18:18]
  wire  _T_1551; // @[CLG.scala 19:18]
  wire  _T_1674; // @[CLG.scala 26:21]
  wire  _T_1675; // @[CLG.scala 26:11]
  wire  _T_1676; // @[CLG.scala 26:31]
  wire  _T_1677; // @[CLG.scala 18:18]
  wire  _T_1678; // @[CLG.scala 19:18]
  wire  _T_1806; // @[CLG.scala 26:21]
  wire  _T_1807; // @[CLG.scala 26:11]
  wire  _T_1808; // @[CLG.scala 26:31]
  wire  _T_1809; // @[CLG.scala 18:18]
  wire  _T_1810; // @[CLG.scala 19:18]
  wire  _T_1943; // @[CLG.scala 26:21]
  wire  _T_1944; // @[CLG.scala 26:11]
  wire  _T_1945; // @[CLG.scala 26:31]
  wire  _T_1946; // @[CLG.scala 18:18]
  wire  _T_1947; // @[CLG.scala 19:18]
  wire  _T_2085; // @[CLG.scala 26:21]
  wire  _T_2086; // @[CLG.scala 26:11]
  wire  _T_2087; // @[CLG.scala 26:31]
  wire  _T_2088; // @[CLG.scala 18:18]
  wire  _T_2089; // @[CLG.scala 19:18]
  wire  _T_2232; // @[CLG.scala 26:21]
  wire  _T_2233; // @[CLG.scala 26:11]
  wire  _T_2234; // @[CLG.scala 26:31]
  wire  _T_2235; // @[CLG.scala 18:18]
  wire  _T_2236; // @[CLG.scala 19:18]
  wire  _T_2384; // @[CLG.scala 26:21]
  wire  _T_2385; // @[CLG.scala 26:11]
  wire  _T_2386; // @[CLG.scala 26:31]
  wire  _T_2387; // @[CLG.scala 18:18]
  wire  _T_2388; // @[CLG.scala 19:18]
  wire  _T_2541; // @[CLG.scala 26:21]
  wire  _T_2542; // @[CLG.scala 26:11]
  wire  _T_2543; // @[CLG.scala 26:31]
  wire  _T_2544; // @[CLG.scala 18:18]
  wire  _T_2545; // @[CLG.scala 19:18]
  wire  _T_2703; // @[CLG.scala 26:21]
  wire  _T_2704; // @[CLG.scala 26:11]
  wire  _T_2705; // @[CLG.scala 26:31]
  wire  _T_2706; // @[CLG.scala 18:18]
  wire  _T_2707; // @[CLG.scala 19:18]
  wire  _T_2870; // @[CLG.scala 26:21]
  wire  _T_2871; // @[CLG.scala 26:11]
  wire  _T_2872; // @[CLG.scala 26:31]
  wire  _T_2873; // @[CLG.scala 18:18]
  wire  _T_2874; // @[CLG.scala 19:18]
  wire  _T_3042; // @[CLG.scala 26:21]
  wire  _T_3043; // @[CLG.scala 26:11]
  wire  _T_3044; // @[CLG.scala 26:31]
  wire  _T_3045; // @[CLG.scala 18:18]
  wire  _T_3046; // @[CLG.scala 19:18]
  wire  _T_3219; // @[CLG.scala 26:21]
  wire  _T_3220; // @[CLG.scala 26:11]
  wire  _T_3221; // @[CLG.scala 26:31]
  wire  _T_3222; // @[CLG.scala 18:18]
  wire  _T_3223; // @[CLG.scala 19:18]
  wire  _T_3401; // @[CLG.scala 26:21]
  wire  _T_3402; // @[CLG.scala 26:11]
  wire  _T_3403; // @[CLG.scala 26:31]
  wire  _T_3404; // @[CLG.scala 18:18]
  wire  _T_3405; // @[CLG.scala 19:18]
  wire  _T_3588; // @[CLG.scala 26:21]
  wire  _T_3589; // @[CLG.scala 26:11]
  wire  _T_3590; // @[CLG.scala 26:31]
  wire  _T_3591; // @[CLG.scala 18:18]
  wire  _T_3592; // @[CLG.scala 19:18]
  wire  _T_3780; // @[CLG.scala 26:21]
  wire  _T_3781; // @[CLG.scala 26:11]
  wire  _T_3782; // @[CLG.scala 26:31]
  wire  _T_3783; // @[CLG.scala 18:18]
  wire  _T_3784; // @[CLG.scala 19:18]
  wire  _T_3977; // @[CLG.scala 26:21]
  wire  _T_3978; // @[CLG.scala 26:11]
  wire  _T_3979; // @[CLG.scala 26:31]
  wire  _T_3980; // @[CLG.scala 18:18]
  wire  _T_3981; // @[CLG.scala 19:18]
  wire  _T_4179; // @[CLG.scala 26:21]
  wire  _T_4180; // @[CLG.scala 26:11]
  wire  _T_4181; // @[CLG.scala 26:31]
  wire  _T_4182; // @[CLG.scala 18:18]
  wire  _T_4183; // @[CLG.scala 19:18]
  wire  _T_4386; // @[CLG.scala 26:21]
  wire  _T_4387; // @[CLG.scala 26:11]
  wire  _T_4388; // @[CLG.scala 26:31]
  wire  _T_4389; // @[CLG.scala 18:18]
  wire  _T_4390; // @[CLG.scala 19:18]
  wire  _T_4598; // @[CLG.scala 26:21]
  wire  _T_4599; // @[CLG.scala 26:11]
  wire  _T_4600; // @[CLG.scala 26:31]
  wire  _T_4601; // @[CLG.scala 18:18]
  wire  _T_4602; // @[CLG.scala 19:18]
  wire  _T_4815; // @[CLG.scala 26:21]
  wire  _T_4816; // @[CLG.scala 26:11]
  wire  _T_4817; // @[CLG.scala 26:31]
  wire  _T_4818; // @[CLG.scala 18:18]
  wire  _T_4819; // @[CLG.scala 19:18]
  wire  _T_5037; // @[CLG.scala 26:21]
  wire  _T_5038; // @[CLG.scala 26:11]
  wire  _T_5039; // @[CLG.scala 26:31]
  wire  _T_5040; // @[CLG.scala 18:18]
  wire  _T_5041; // @[CLG.scala 19:18]
  wire  _T_5264; // @[CLG.scala 26:21]
  wire  _T_5265; // @[CLG.scala 26:11]
  wire  _T_5266; // @[CLG.scala 26:31]
  wire  _T_5267; // @[CLG.scala 18:18]
  wire  _T_5268; // @[CLG.scala 19:18]
  wire  _T_5496; // @[CLG.scala 26:21]
  wire  _T_5497; // @[CLG.scala 26:11]
  wire  _T_5498; // @[CLG.scala 26:31]
  wire  _T_5499; // @[CLG.scala 18:18]
  wire  _T_5500; // @[CLG.scala 19:18]
  wire  _T_5733; // @[CLG.scala 26:21]
  wire  _T_5734; // @[CLG.scala 26:11]
  wire  _T_5735; // @[CLG.scala 26:31]
  wire  _T_5736; // @[CLG.scala 18:18]
  wire  _T_5737; // @[CLG.scala 19:18]
  wire  _T_5975; // @[CLG.scala 26:21]
  wire  _T_5976; // @[CLG.scala 26:11]
  wire  _T_5977; // @[CLG.scala 26:31]
  wire  _T_5978; // @[CLG.scala 18:18]
  wire  _T_5979; // @[CLG.scala 19:18]
  wire  _T_6222; // @[CLG.scala 26:21]
  wire  _T_6223; // @[CLG.scala 26:11]
  wire  _T_6224; // @[CLG.scala 26:31]
  wire  _T_6225; // @[CLG.scala 18:18]
  wire  _T_6226; // @[CLG.scala 19:18]
  wire  _T_6474; // @[CLG.scala 26:21]
  wire  _T_6475; // @[CLG.scala 26:11]
  wire  _T_6476; // @[CLG.scala 26:31]
  wire  _T_6477; // @[CLG.scala 18:18]
  wire  _T_6478; // @[CLG.scala 19:18]
  wire  _T_6731; // @[CLG.scala 26:21]
  wire  _T_6732; // @[CLG.scala 26:11]
  wire  _T_6733; // @[CLG.scala 26:31]
  wire  _T_6734; // @[CLG.scala 18:18]
  wire  _T_6735; // @[CLG.scala 19:18]
  wire  _T_6993; // @[CLG.scala 26:21]
  wire  _T_6994; // @[CLG.scala 26:11]
  wire  _T_6995; // @[CLG.scala 26:31]
  wire  _T_6996; // @[CLG.scala 18:18]
  wire  _T_6997; // @[CLG.scala 19:18]
  wire  _T_7260; // @[CLG.scala 26:21]
  wire  _T_7261; // @[CLG.scala 26:11]
  wire  _T_7262; // @[CLG.scala 26:31]
  wire  _T_7263; // @[CLG.scala 18:18]
  wire  _T_7264; // @[CLG.scala 19:18]
  wire  _T_7532; // @[CLG.scala 26:21]
  wire  _T_7533; // @[CLG.scala 26:11]
  wire  _T_7534; // @[CLG.scala 26:31]
  wire  _T_7535; // @[CLG.scala 18:18]
  wire  _T_7536; // @[CLG.scala 19:18]
  wire  _T_7809; // @[CLG.scala 26:21]
  wire  _T_7810; // @[CLG.scala 26:11]
  wire  _T_7811; // @[CLG.scala 26:31]
  wire  _T_7812; // @[CLG.scala 18:18]
  wire  _T_7813; // @[CLG.scala 19:18]
  wire  _T_8091; // @[CLG.scala 26:21]
  wire  _T_8092; // @[CLG.scala 26:11]
  wire  _T_8093; // @[CLG.scala 26:31]
  wire  _T_8094; // @[CLG.scala 18:18]
  wire  _T_8095; // @[CLG.scala 19:18]
  wire  _T_8378; // @[CLG.scala 26:21]
  wire  _T_8379; // @[CLG.scala 26:11]
  wire  _T_8380; // @[CLG.scala 26:31]
  wire  _T_8381; // @[CLG.scala 18:18]
  wire  _T_8382; // @[CLG.scala 19:18]
  wire  _T_8670; // @[CLG.scala 26:21]
  wire  _T_8671; // @[CLG.scala 26:11]
  wire  _T_8672; // @[CLG.scala 26:31]
  wire  _T_8673; // @[CLG.scala 18:18]
  wire  _T_8674; // @[CLG.scala 19:18]
  wire  _T_8967; // @[CLG.scala 26:21]
  wire  _T_8968; // @[CLG.scala 26:11]
  wire  _T_8969; // @[CLG.scala 26:31]
  wire  _T_8970; // @[CLG.scala 18:18]
  wire  _T_8971; // @[CLG.scala 19:18]
  wire  _T_9269; // @[CLG.scala 26:21]
  wire  _T_9270; // @[CLG.scala 26:11]
  wire  _T_9271; // @[CLG.scala 26:31]
  wire  _T_9272; // @[CLG.scala 18:18]
  wire  _T_9273; // @[CLG.scala 19:18]
  wire  _T_9576; // @[CLG.scala 26:21]
  wire  _T_9577; // @[CLG.scala 26:11]
  wire  _T_9578; // @[CLG.scala 26:31]
  wire  _T_9579; // @[CLG.scala 18:18]
  wire  _T_9580; // @[CLG.scala 19:18]
  wire  _T_9888; // @[CLG.scala 26:21]
  wire  _T_9889; // @[CLG.scala 26:11]
  wire  _T_9890; // @[CLG.scala 26:31]
  wire  _T_9891; // @[CLG.scala 18:18]
  wire  _T_9892; // @[CLG.scala 19:18]
  wire  _T_10205; // @[CLG.scala 26:21]
  wire  _T_10206; // @[CLG.scala 26:11]
  wire  _T_10207; // @[CLG.scala 26:31]
  wire  _T_10208; // @[CLG.scala 41:22]
  wire  c_bit_0; // @[CLG.scala 41:12]
  wire  _T_10209; // @[CLG.scala 41:22]
  wire  c_bit_1; // @[CLG.scala 41:12]
  wire  _T_10210; // @[CLG.scala 41:22]
  wire  c_bit_2; // @[CLG.scala 41:12]
  wire  _T_10211; // @[CLG.scala 41:22]
  wire  c_bit_3; // @[CLG.scala 41:12]
  wire  _T_10212; // @[CLG.scala 41:22]
  wire  c_bit_4; // @[CLG.scala 41:12]
  wire  _T_10213; // @[CLG.scala 41:22]
  wire  c_bit_5; // @[CLG.scala 41:12]
  wire  _T_10214; // @[CLG.scala 41:22]
  wire  c_bit_6; // @[CLG.scala 41:12]
  wire  _T_10215; // @[CLG.scala 41:22]
  wire  c_bit_7; // @[CLG.scala 41:12]
  wire  _T_10216; // @[CLG.scala 41:22]
  wire  c_bit_8; // @[CLG.scala 41:12]
  wire  _T_10217; // @[CLG.scala 41:22]
  wire  c_bit_9; // @[CLG.scala 41:12]
  wire  _T_10218; // @[CLG.scala 41:22]
  wire  c_bit_10; // @[CLG.scala 41:12]
  wire  _T_10219; // @[CLG.scala 41:22]
  wire  c_bit_11; // @[CLG.scala 41:12]
  wire  _T_10220; // @[CLG.scala 41:22]
  wire  c_bit_12; // @[CLG.scala 41:12]
  wire  _T_10221; // @[CLG.scala 41:22]
  wire  c_bit_13; // @[CLG.scala 41:12]
  wire  _T_10222; // @[CLG.scala 41:22]
  wire  c_bit_14; // @[CLG.scala 41:12]
  wire  _T_10223; // @[CLG.scala 41:22]
  wire  c_bit_15; // @[CLG.scala 41:12]
  wire  _T_10224; // @[CLG.scala 41:22]
  wire  c_bit_16; // @[CLG.scala 41:12]
  wire  _T_10225; // @[CLG.scala 41:22]
  wire  c_bit_17; // @[CLG.scala 41:12]
  wire  _T_10226; // @[CLG.scala 41:22]
  wire  c_bit_18; // @[CLG.scala 41:12]
  wire  _T_10227; // @[CLG.scala 41:22]
  wire  c_bit_19; // @[CLG.scala 41:12]
  wire  _T_10228; // @[CLG.scala 41:22]
  wire  c_bit_20; // @[CLG.scala 41:12]
  wire  _T_10229; // @[CLG.scala 41:22]
  wire  c_bit_21; // @[CLG.scala 41:12]
  wire  _T_10230; // @[CLG.scala 41:22]
  wire  c_bit_22; // @[CLG.scala 41:12]
  wire  _T_10231; // @[CLG.scala 41:22]
  wire  c_bit_23; // @[CLG.scala 41:12]
  wire  _T_10232; // @[CLG.scala 41:22]
  wire  c_bit_24; // @[CLG.scala 41:12]
  wire  _T_10233; // @[CLG.scala 41:22]
  wire  c_bit_25; // @[CLG.scala 41:12]
  wire  _T_10234; // @[CLG.scala 41:22]
  wire  c_bit_26; // @[CLG.scala 41:12]
  wire  _T_10235; // @[CLG.scala 41:22]
  wire  c_bit_27; // @[CLG.scala 41:12]
  wire  _T_10236; // @[CLG.scala 41:22]
  wire  c_bit_28; // @[CLG.scala 41:12]
  wire  _T_10237; // @[CLG.scala 41:22]
  wire  c_bit_29; // @[CLG.scala 41:12]
  wire  _T_10238; // @[CLG.scala 41:22]
  wire  c_bit_30; // @[CLG.scala 41:12]
  wire  _T_10239; // @[CLG.scala 41:22]
  wire  c_bit_31; // @[CLG.scala 41:12]
  wire  _T_10240; // @[CLG.scala 41:22]
  wire  c_bit_32; // @[CLG.scala 41:12]
  wire  _T_10241; // @[CLG.scala 41:22]
  wire  c_bit_33; // @[CLG.scala 41:12]
  wire  _T_10242; // @[CLG.scala 41:22]
  wire  c_bit_34; // @[CLG.scala 41:12]
  wire  _T_10243; // @[CLG.scala 41:22]
  wire  c_bit_35; // @[CLG.scala 41:12]
  wire  _T_10244; // @[CLG.scala 41:22]
  wire  c_bit_36; // @[CLG.scala 41:12]
  wire  _T_10245; // @[CLG.scala 41:22]
  wire  c_bit_37; // @[CLG.scala 41:12]
  wire  _T_10246; // @[CLG.scala 41:22]
  wire  c_bit_38; // @[CLG.scala 41:12]
  wire  _T_10247; // @[CLG.scala 41:22]
  wire  c_bit_39; // @[CLG.scala 41:12]
  wire  _T_10248; // @[CLG.scala 41:22]
  wire  c_bit_40; // @[CLG.scala 41:12]
  wire  _T_10249; // @[CLG.scala 41:22]
  wire  c_bit_41; // @[CLG.scala 41:12]
  wire  _T_10250; // @[CLG.scala 41:22]
  wire  c_bit_42; // @[CLG.scala 41:12]
  wire  _T_10251; // @[CLG.scala 41:22]
  wire  c_bit_43; // @[CLG.scala 41:12]
  wire  _T_10252; // @[CLG.scala 41:22]
  wire  c_bit_44; // @[CLG.scala 41:12]
  wire  _T_10253; // @[CLG.scala 41:22]
  wire  c_bit_45; // @[CLG.scala 41:12]
  wire  _T_10254; // @[CLG.scala 41:22]
  wire  c_bit_46; // @[CLG.scala 41:12]
  wire  _T_10255; // @[CLG.scala 41:22]
  wire  c_bit_47; // @[CLG.scala 41:12]
  wire  _T_10256; // @[CLG.scala 41:22]
  wire  c_bit_48; // @[CLG.scala 41:12]
  wire  _T_10257; // @[CLG.scala 41:22]
  wire  c_bit_49; // @[CLG.scala 41:12]
  wire  _T_10258; // @[CLG.scala 41:22]
  wire  c_bit_50; // @[CLG.scala 41:12]
  wire  _T_10259; // @[CLG.scala 41:22]
  wire  c_bit_51; // @[CLG.scala 41:12]
  wire  _T_10260; // @[CLG.scala 41:22]
  wire  c_bit_52; // @[CLG.scala 41:12]
  wire  _T_10261; // @[CLG.scala 41:22]
  wire  c_bit_53; // @[CLG.scala 41:12]
  wire  _T_10262; // @[CLG.scala 41:22]
  wire  c_bit_54; // @[CLG.scala 41:12]
  wire  _T_10263; // @[CLG.scala 41:22]
  wire  c_bit_55; // @[CLG.scala 41:12]
  wire  _T_10264; // @[CLG.scala 41:22]
  wire  c_bit_56; // @[CLG.scala 41:12]
  wire  _T_10265; // @[CLG.scala 41:22]
  wire  c_bit_57; // @[CLG.scala 41:12]
  wire  _T_10266; // @[CLG.scala 41:22]
  wire  c_bit_58; // @[CLG.scala 41:12]
  wire  _T_10267; // @[CLG.scala 41:22]
  wire  c_bit_59; // @[CLG.scala 41:12]
  wire  _T_10268; // @[CLG.scala 41:22]
  wire  c_bit_60; // @[CLG.scala 41:12]
  wire  _T_10269; // @[CLG.scala 41:22]
  wire  c_bit_61; // @[CLG.scala 41:12]
  wire  _T_10270; // @[CLG.scala 41:22]
  wire  c_bit_62; // @[CLG.scala 41:12]
  wire  _T_10271; // @[CLG.scala 41:22]
  wire  c_bit_63; // @[CLG.scala 41:12]
  wire [7:0] _T_10279; // @[CLG.scala 43:32]
  wire [15:0] _T_10287; // @[CLG.scala 43:32]
  wire [7:0] _T_10294; // @[CLG.scala 43:32]
  wire [31:0] _T_10303; // @[CLG.scala 43:32]
  wire [7:0] _T_10310; // @[CLG.scala 43:32]
  wire [15:0] _T_10318; // @[CLG.scala 43:32]
  wire [7:0] _T_10325; // @[CLG.scala 43:32]
  wire [31:0] _T_10334; // @[CLG.scala 43:32]
  assign _T = io_g[0]; // @[CLG.scala 18:18]
  assign _T_1 = io_a[0]; // @[CLG.scala 19:18]
  assign _T_2 = io_g[1]; // @[CLG.scala 18:18]
  assign _T_3 = io_a[1]; // @[CLG.scala 19:18]
  assign _T_6 = _T & _T_3; // @[CLG.scala 26:21]
  assign _T_7 = _T_2 | _T_6; // @[CLG.scala 26:11]
  assign _T_8 = _T_3 & _T_1; // @[CLG.scala 26:31]
  assign _T_9 = io_g[2]; // @[CLG.scala 18:18]
  assign _T_10 = io_a[2]; // @[CLG.scala 19:18]
  assign _T_18 = _T_7 & _T_10; // @[CLG.scala 26:21]
  assign _T_19 = _T_9 | _T_18; // @[CLG.scala 26:11]
  assign _T_20 = _T_10 & _T_8; // @[CLG.scala 26:31]
  assign _T_21 = io_g[3]; // @[CLG.scala 18:18]
  assign _T_22 = io_a[3]; // @[CLG.scala 19:18]
  assign _T_35 = _T_19 & _T_22; // @[CLG.scala 26:21]
  assign _T_36 = _T_21 | _T_35; // @[CLG.scala 26:11]
  assign _T_37 = _T_22 & _T_20; // @[CLG.scala 26:31]
  assign _T_38 = io_g[4]; // @[CLG.scala 18:18]
  assign _T_39 = io_a[4]; // @[CLG.scala 19:18]
  assign _T_57 = _T_36 & _T_39; // @[CLG.scala 26:21]
  assign _T_58 = _T_38 | _T_57; // @[CLG.scala 26:11]
  assign _T_59 = _T_39 & _T_37; // @[CLG.scala 26:31]
  assign _T_60 = io_g[5]; // @[CLG.scala 18:18]
  assign _T_61 = io_a[5]; // @[CLG.scala 19:18]
  assign _T_84 = _T_58 & _T_61; // @[CLG.scala 26:21]
  assign _T_85 = _T_60 | _T_84; // @[CLG.scala 26:11]
  assign _T_86 = _T_61 & _T_59; // @[CLG.scala 26:31]
  assign _T_87 = io_g[6]; // @[CLG.scala 18:18]
  assign _T_88 = io_a[6]; // @[CLG.scala 19:18]
  assign _T_116 = _T_85 & _T_88; // @[CLG.scala 26:21]
  assign _T_117 = _T_87 | _T_116; // @[CLG.scala 26:11]
  assign _T_118 = _T_88 & _T_86; // @[CLG.scala 26:31]
  assign _T_119 = io_g[7]; // @[CLG.scala 18:18]
  assign _T_120 = io_a[7]; // @[CLG.scala 19:18]
  assign _T_153 = _T_117 & _T_120; // @[CLG.scala 26:21]
  assign _T_154 = _T_119 | _T_153; // @[CLG.scala 26:11]
  assign _T_155 = _T_120 & _T_118; // @[CLG.scala 26:31]
  assign _T_156 = io_g[8]; // @[CLG.scala 18:18]
  assign _T_157 = io_a[8]; // @[CLG.scala 19:18]
  assign _T_195 = _T_154 & _T_157; // @[CLG.scala 26:21]
  assign _T_196 = _T_156 | _T_195; // @[CLG.scala 26:11]
  assign _T_197 = _T_157 & _T_155; // @[CLG.scala 26:31]
  assign _T_198 = io_g[9]; // @[CLG.scala 18:18]
  assign _T_199 = io_a[9]; // @[CLG.scala 19:18]
  assign _T_242 = _T_196 & _T_199; // @[CLG.scala 26:21]
  assign _T_243 = _T_198 | _T_242; // @[CLG.scala 26:11]
  assign _T_244 = _T_199 & _T_197; // @[CLG.scala 26:31]
  assign _T_245 = io_g[10]; // @[CLG.scala 18:18]
  assign _T_246 = io_a[10]; // @[CLG.scala 19:18]
  assign _T_294 = _T_243 & _T_246; // @[CLG.scala 26:21]
  assign _T_295 = _T_245 | _T_294; // @[CLG.scala 26:11]
  assign _T_296 = _T_246 & _T_244; // @[CLG.scala 26:31]
  assign _T_297 = io_g[11]; // @[CLG.scala 18:18]
  assign _T_298 = io_a[11]; // @[CLG.scala 19:18]
  assign _T_351 = _T_295 & _T_298; // @[CLG.scala 26:21]
  assign _T_352 = _T_297 | _T_351; // @[CLG.scala 26:11]
  assign _T_353 = _T_298 & _T_296; // @[CLG.scala 26:31]
  assign _T_354 = io_g[12]; // @[CLG.scala 18:18]
  assign _T_355 = io_a[12]; // @[CLG.scala 19:18]
  assign _T_413 = _T_352 & _T_355; // @[CLG.scala 26:21]
  assign _T_414 = _T_354 | _T_413; // @[CLG.scala 26:11]
  assign _T_415 = _T_355 & _T_353; // @[CLG.scala 26:31]
  assign _T_416 = io_g[13]; // @[CLG.scala 18:18]
  assign _T_417 = io_a[13]; // @[CLG.scala 19:18]
  assign _T_480 = _T_414 & _T_417; // @[CLG.scala 26:21]
  assign _T_481 = _T_416 | _T_480; // @[CLG.scala 26:11]
  assign _T_482 = _T_417 & _T_415; // @[CLG.scala 26:31]
  assign _T_483 = io_g[14]; // @[CLG.scala 18:18]
  assign _T_484 = io_a[14]; // @[CLG.scala 19:18]
  assign _T_552 = _T_481 & _T_484; // @[CLG.scala 26:21]
  assign _T_553 = _T_483 | _T_552; // @[CLG.scala 26:11]
  assign _T_554 = _T_484 & _T_482; // @[CLG.scala 26:31]
  assign _T_555 = io_g[15]; // @[CLG.scala 18:18]
  assign _T_556 = io_a[15]; // @[CLG.scala 19:18]
  assign _T_629 = _T_553 & _T_556; // @[CLG.scala 26:21]
  assign _T_630 = _T_555 | _T_629; // @[CLG.scala 26:11]
  assign _T_631 = _T_556 & _T_554; // @[CLG.scala 26:31]
  assign _T_632 = io_g[16]; // @[CLG.scala 18:18]
  assign _T_633 = io_a[16]; // @[CLG.scala 19:18]
  assign _T_711 = _T_630 & _T_633; // @[CLG.scala 26:21]
  assign _T_712 = _T_632 | _T_711; // @[CLG.scala 26:11]
  assign _T_713 = _T_633 & _T_631; // @[CLG.scala 26:31]
  assign _T_714 = io_g[17]; // @[CLG.scala 18:18]
  assign _T_715 = io_a[17]; // @[CLG.scala 19:18]
  assign _T_798 = _T_712 & _T_715; // @[CLG.scala 26:21]
  assign _T_799 = _T_714 | _T_798; // @[CLG.scala 26:11]
  assign _T_800 = _T_715 & _T_713; // @[CLG.scala 26:31]
  assign _T_801 = io_g[18]; // @[CLG.scala 18:18]
  assign _T_802 = io_a[18]; // @[CLG.scala 19:18]
  assign _T_890 = _T_799 & _T_802; // @[CLG.scala 26:21]
  assign _T_891 = _T_801 | _T_890; // @[CLG.scala 26:11]
  assign _T_892 = _T_802 & _T_800; // @[CLG.scala 26:31]
  assign _T_893 = io_g[19]; // @[CLG.scala 18:18]
  assign _T_894 = io_a[19]; // @[CLG.scala 19:18]
  assign _T_987 = _T_891 & _T_894; // @[CLG.scala 26:21]
  assign _T_988 = _T_893 | _T_987; // @[CLG.scala 26:11]
  assign _T_989 = _T_894 & _T_892; // @[CLG.scala 26:31]
  assign _T_990 = io_g[20]; // @[CLG.scala 18:18]
  assign _T_991 = io_a[20]; // @[CLG.scala 19:18]
  assign _T_1089 = _T_988 & _T_991; // @[CLG.scala 26:21]
  assign _T_1090 = _T_990 | _T_1089; // @[CLG.scala 26:11]
  assign _T_1091 = _T_991 & _T_989; // @[CLG.scala 26:31]
  assign _T_1092 = io_g[21]; // @[CLG.scala 18:18]
  assign _T_1093 = io_a[21]; // @[CLG.scala 19:18]
  assign _T_1196 = _T_1090 & _T_1093; // @[CLG.scala 26:21]
  assign _T_1197 = _T_1092 | _T_1196; // @[CLG.scala 26:11]
  assign _T_1198 = _T_1093 & _T_1091; // @[CLG.scala 26:31]
  assign _T_1199 = io_g[22]; // @[CLG.scala 18:18]
  assign _T_1200 = io_a[22]; // @[CLG.scala 19:18]
  assign _T_1308 = _T_1197 & _T_1200; // @[CLG.scala 26:21]
  assign _T_1309 = _T_1199 | _T_1308; // @[CLG.scala 26:11]
  assign _T_1310 = _T_1200 & _T_1198; // @[CLG.scala 26:31]
  assign _T_1311 = io_g[23]; // @[CLG.scala 18:18]
  assign _T_1312 = io_a[23]; // @[CLG.scala 19:18]
  assign _T_1425 = _T_1309 & _T_1312; // @[CLG.scala 26:21]
  assign _T_1426 = _T_1311 | _T_1425; // @[CLG.scala 26:11]
  assign _T_1427 = _T_1312 & _T_1310; // @[CLG.scala 26:31]
  assign _T_1428 = io_g[24]; // @[CLG.scala 18:18]
  assign _T_1429 = io_a[24]; // @[CLG.scala 19:18]
  assign _T_1547 = _T_1426 & _T_1429; // @[CLG.scala 26:21]
  assign _T_1548 = _T_1428 | _T_1547; // @[CLG.scala 26:11]
  assign _T_1549 = _T_1429 & _T_1427; // @[CLG.scala 26:31]
  assign _T_1550 = io_g[25]; // @[CLG.scala 18:18]
  assign _T_1551 = io_a[25]; // @[CLG.scala 19:18]
  assign _T_1674 = _T_1548 & _T_1551; // @[CLG.scala 26:21]
  assign _T_1675 = _T_1550 | _T_1674; // @[CLG.scala 26:11]
  assign _T_1676 = _T_1551 & _T_1549; // @[CLG.scala 26:31]
  assign _T_1677 = io_g[26]; // @[CLG.scala 18:18]
  assign _T_1678 = io_a[26]; // @[CLG.scala 19:18]
  assign _T_1806 = _T_1675 & _T_1678; // @[CLG.scala 26:21]
  assign _T_1807 = _T_1677 | _T_1806; // @[CLG.scala 26:11]
  assign _T_1808 = _T_1678 & _T_1676; // @[CLG.scala 26:31]
  assign _T_1809 = io_g[27]; // @[CLG.scala 18:18]
  assign _T_1810 = io_a[27]; // @[CLG.scala 19:18]
  assign _T_1943 = _T_1807 & _T_1810; // @[CLG.scala 26:21]
  assign _T_1944 = _T_1809 | _T_1943; // @[CLG.scala 26:11]
  assign _T_1945 = _T_1810 & _T_1808; // @[CLG.scala 26:31]
  assign _T_1946 = io_g[28]; // @[CLG.scala 18:18]
  assign _T_1947 = io_a[28]; // @[CLG.scala 19:18]
  assign _T_2085 = _T_1944 & _T_1947; // @[CLG.scala 26:21]
  assign _T_2086 = _T_1946 | _T_2085; // @[CLG.scala 26:11]
  assign _T_2087 = _T_1947 & _T_1945; // @[CLG.scala 26:31]
  assign _T_2088 = io_g[29]; // @[CLG.scala 18:18]
  assign _T_2089 = io_a[29]; // @[CLG.scala 19:18]
  assign _T_2232 = _T_2086 & _T_2089; // @[CLG.scala 26:21]
  assign _T_2233 = _T_2088 | _T_2232; // @[CLG.scala 26:11]
  assign _T_2234 = _T_2089 & _T_2087; // @[CLG.scala 26:31]
  assign _T_2235 = io_g[30]; // @[CLG.scala 18:18]
  assign _T_2236 = io_a[30]; // @[CLG.scala 19:18]
  assign _T_2384 = _T_2233 & _T_2236; // @[CLG.scala 26:21]
  assign _T_2385 = _T_2235 | _T_2384; // @[CLG.scala 26:11]
  assign _T_2386 = _T_2236 & _T_2234; // @[CLG.scala 26:31]
  assign _T_2387 = io_g[31]; // @[CLG.scala 18:18]
  assign _T_2388 = io_a[31]; // @[CLG.scala 19:18]
  assign _T_2541 = _T_2385 & _T_2388; // @[CLG.scala 26:21]
  assign _T_2542 = _T_2387 | _T_2541; // @[CLG.scala 26:11]
  assign _T_2543 = _T_2388 & _T_2386; // @[CLG.scala 26:31]
  assign _T_2544 = io_g[32]; // @[CLG.scala 18:18]
  assign _T_2545 = io_a[32]; // @[CLG.scala 19:18]
  assign _T_2703 = _T_2542 & _T_2545; // @[CLG.scala 26:21]
  assign _T_2704 = _T_2544 | _T_2703; // @[CLG.scala 26:11]
  assign _T_2705 = _T_2545 & _T_2543; // @[CLG.scala 26:31]
  assign _T_2706 = io_g[33]; // @[CLG.scala 18:18]
  assign _T_2707 = io_a[33]; // @[CLG.scala 19:18]
  assign _T_2870 = _T_2704 & _T_2707; // @[CLG.scala 26:21]
  assign _T_2871 = _T_2706 | _T_2870; // @[CLG.scala 26:11]
  assign _T_2872 = _T_2707 & _T_2705; // @[CLG.scala 26:31]
  assign _T_2873 = io_g[34]; // @[CLG.scala 18:18]
  assign _T_2874 = io_a[34]; // @[CLG.scala 19:18]
  assign _T_3042 = _T_2871 & _T_2874; // @[CLG.scala 26:21]
  assign _T_3043 = _T_2873 | _T_3042; // @[CLG.scala 26:11]
  assign _T_3044 = _T_2874 & _T_2872; // @[CLG.scala 26:31]
  assign _T_3045 = io_g[35]; // @[CLG.scala 18:18]
  assign _T_3046 = io_a[35]; // @[CLG.scala 19:18]
  assign _T_3219 = _T_3043 & _T_3046; // @[CLG.scala 26:21]
  assign _T_3220 = _T_3045 | _T_3219; // @[CLG.scala 26:11]
  assign _T_3221 = _T_3046 & _T_3044; // @[CLG.scala 26:31]
  assign _T_3222 = io_g[36]; // @[CLG.scala 18:18]
  assign _T_3223 = io_a[36]; // @[CLG.scala 19:18]
  assign _T_3401 = _T_3220 & _T_3223; // @[CLG.scala 26:21]
  assign _T_3402 = _T_3222 | _T_3401; // @[CLG.scala 26:11]
  assign _T_3403 = _T_3223 & _T_3221; // @[CLG.scala 26:31]
  assign _T_3404 = io_g[37]; // @[CLG.scala 18:18]
  assign _T_3405 = io_a[37]; // @[CLG.scala 19:18]
  assign _T_3588 = _T_3402 & _T_3405; // @[CLG.scala 26:21]
  assign _T_3589 = _T_3404 | _T_3588; // @[CLG.scala 26:11]
  assign _T_3590 = _T_3405 & _T_3403; // @[CLG.scala 26:31]
  assign _T_3591 = io_g[38]; // @[CLG.scala 18:18]
  assign _T_3592 = io_a[38]; // @[CLG.scala 19:18]
  assign _T_3780 = _T_3589 & _T_3592; // @[CLG.scala 26:21]
  assign _T_3781 = _T_3591 | _T_3780; // @[CLG.scala 26:11]
  assign _T_3782 = _T_3592 & _T_3590; // @[CLG.scala 26:31]
  assign _T_3783 = io_g[39]; // @[CLG.scala 18:18]
  assign _T_3784 = io_a[39]; // @[CLG.scala 19:18]
  assign _T_3977 = _T_3781 & _T_3784; // @[CLG.scala 26:21]
  assign _T_3978 = _T_3783 | _T_3977; // @[CLG.scala 26:11]
  assign _T_3979 = _T_3784 & _T_3782; // @[CLG.scala 26:31]
  assign _T_3980 = io_g[40]; // @[CLG.scala 18:18]
  assign _T_3981 = io_a[40]; // @[CLG.scala 19:18]
  assign _T_4179 = _T_3978 & _T_3981; // @[CLG.scala 26:21]
  assign _T_4180 = _T_3980 | _T_4179; // @[CLG.scala 26:11]
  assign _T_4181 = _T_3981 & _T_3979; // @[CLG.scala 26:31]
  assign _T_4182 = io_g[41]; // @[CLG.scala 18:18]
  assign _T_4183 = io_a[41]; // @[CLG.scala 19:18]
  assign _T_4386 = _T_4180 & _T_4183; // @[CLG.scala 26:21]
  assign _T_4387 = _T_4182 | _T_4386; // @[CLG.scala 26:11]
  assign _T_4388 = _T_4183 & _T_4181; // @[CLG.scala 26:31]
  assign _T_4389 = io_g[42]; // @[CLG.scala 18:18]
  assign _T_4390 = io_a[42]; // @[CLG.scala 19:18]
  assign _T_4598 = _T_4387 & _T_4390; // @[CLG.scala 26:21]
  assign _T_4599 = _T_4389 | _T_4598; // @[CLG.scala 26:11]
  assign _T_4600 = _T_4390 & _T_4388; // @[CLG.scala 26:31]
  assign _T_4601 = io_g[43]; // @[CLG.scala 18:18]
  assign _T_4602 = io_a[43]; // @[CLG.scala 19:18]
  assign _T_4815 = _T_4599 & _T_4602; // @[CLG.scala 26:21]
  assign _T_4816 = _T_4601 | _T_4815; // @[CLG.scala 26:11]
  assign _T_4817 = _T_4602 & _T_4600; // @[CLG.scala 26:31]
  assign _T_4818 = io_g[44]; // @[CLG.scala 18:18]
  assign _T_4819 = io_a[44]; // @[CLG.scala 19:18]
  assign _T_5037 = _T_4816 & _T_4819; // @[CLG.scala 26:21]
  assign _T_5038 = _T_4818 | _T_5037; // @[CLG.scala 26:11]
  assign _T_5039 = _T_4819 & _T_4817; // @[CLG.scala 26:31]
  assign _T_5040 = io_g[45]; // @[CLG.scala 18:18]
  assign _T_5041 = io_a[45]; // @[CLG.scala 19:18]
  assign _T_5264 = _T_5038 & _T_5041; // @[CLG.scala 26:21]
  assign _T_5265 = _T_5040 | _T_5264; // @[CLG.scala 26:11]
  assign _T_5266 = _T_5041 & _T_5039; // @[CLG.scala 26:31]
  assign _T_5267 = io_g[46]; // @[CLG.scala 18:18]
  assign _T_5268 = io_a[46]; // @[CLG.scala 19:18]
  assign _T_5496 = _T_5265 & _T_5268; // @[CLG.scala 26:21]
  assign _T_5497 = _T_5267 | _T_5496; // @[CLG.scala 26:11]
  assign _T_5498 = _T_5268 & _T_5266; // @[CLG.scala 26:31]
  assign _T_5499 = io_g[47]; // @[CLG.scala 18:18]
  assign _T_5500 = io_a[47]; // @[CLG.scala 19:18]
  assign _T_5733 = _T_5497 & _T_5500; // @[CLG.scala 26:21]
  assign _T_5734 = _T_5499 | _T_5733; // @[CLG.scala 26:11]
  assign _T_5735 = _T_5500 & _T_5498; // @[CLG.scala 26:31]
  assign _T_5736 = io_g[48]; // @[CLG.scala 18:18]
  assign _T_5737 = io_a[48]; // @[CLG.scala 19:18]
  assign _T_5975 = _T_5734 & _T_5737; // @[CLG.scala 26:21]
  assign _T_5976 = _T_5736 | _T_5975; // @[CLG.scala 26:11]
  assign _T_5977 = _T_5737 & _T_5735; // @[CLG.scala 26:31]
  assign _T_5978 = io_g[49]; // @[CLG.scala 18:18]
  assign _T_5979 = io_a[49]; // @[CLG.scala 19:18]
  assign _T_6222 = _T_5976 & _T_5979; // @[CLG.scala 26:21]
  assign _T_6223 = _T_5978 | _T_6222; // @[CLG.scala 26:11]
  assign _T_6224 = _T_5979 & _T_5977; // @[CLG.scala 26:31]
  assign _T_6225 = io_g[50]; // @[CLG.scala 18:18]
  assign _T_6226 = io_a[50]; // @[CLG.scala 19:18]
  assign _T_6474 = _T_6223 & _T_6226; // @[CLG.scala 26:21]
  assign _T_6475 = _T_6225 | _T_6474; // @[CLG.scala 26:11]
  assign _T_6476 = _T_6226 & _T_6224; // @[CLG.scala 26:31]
  assign _T_6477 = io_g[51]; // @[CLG.scala 18:18]
  assign _T_6478 = io_a[51]; // @[CLG.scala 19:18]
  assign _T_6731 = _T_6475 & _T_6478; // @[CLG.scala 26:21]
  assign _T_6732 = _T_6477 | _T_6731; // @[CLG.scala 26:11]
  assign _T_6733 = _T_6478 & _T_6476; // @[CLG.scala 26:31]
  assign _T_6734 = io_g[52]; // @[CLG.scala 18:18]
  assign _T_6735 = io_a[52]; // @[CLG.scala 19:18]
  assign _T_6993 = _T_6732 & _T_6735; // @[CLG.scala 26:21]
  assign _T_6994 = _T_6734 | _T_6993; // @[CLG.scala 26:11]
  assign _T_6995 = _T_6735 & _T_6733; // @[CLG.scala 26:31]
  assign _T_6996 = io_g[53]; // @[CLG.scala 18:18]
  assign _T_6997 = io_a[53]; // @[CLG.scala 19:18]
  assign _T_7260 = _T_6994 & _T_6997; // @[CLG.scala 26:21]
  assign _T_7261 = _T_6996 | _T_7260; // @[CLG.scala 26:11]
  assign _T_7262 = _T_6997 & _T_6995; // @[CLG.scala 26:31]
  assign _T_7263 = io_g[54]; // @[CLG.scala 18:18]
  assign _T_7264 = io_a[54]; // @[CLG.scala 19:18]
  assign _T_7532 = _T_7261 & _T_7264; // @[CLG.scala 26:21]
  assign _T_7533 = _T_7263 | _T_7532; // @[CLG.scala 26:11]
  assign _T_7534 = _T_7264 & _T_7262; // @[CLG.scala 26:31]
  assign _T_7535 = io_g[55]; // @[CLG.scala 18:18]
  assign _T_7536 = io_a[55]; // @[CLG.scala 19:18]
  assign _T_7809 = _T_7533 & _T_7536; // @[CLG.scala 26:21]
  assign _T_7810 = _T_7535 | _T_7809; // @[CLG.scala 26:11]
  assign _T_7811 = _T_7536 & _T_7534; // @[CLG.scala 26:31]
  assign _T_7812 = io_g[56]; // @[CLG.scala 18:18]
  assign _T_7813 = io_a[56]; // @[CLG.scala 19:18]
  assign _T_8091 = _T_7810 & _T_7813; // @[CLG.scala 26:21]
  assign _T_8092 = _T_7812 | _T_8091; // @[CLG.scala 26:11]
  assign _T_8093 = _T_7813 & _T_7811; // @[CLG.scala 26:31]
  assign _T_8094 = io_g[57]; // @[CLG.scala 18:18]
  assign _T_8095 = io_a[57]; // @[CLG.scala 19:18]
  assign _T_8378 = _T_8092 & _T_8095; // @[CLG.scala 26:21]
  assign _T_8379 = _T_8094 | _T_8378; // @[CLG.scala 26:11]
  assign _T_8380 = _T_8095 & _T_8093; // @[CLG.scala 26:31]
  assign _T_8381 = io_g[58]; // @[CLG.scala 18:18]
  assign _T_8382 = io_a[58]; // @[CLG.scala 19:18]
  assign _T_8670 = _T_8379 & _T_8382; // @[CLG.scala 26:21]
  assign _T_8671 = _T_8381 | _T_8670; // @[CLG.scala 26:11]
  assign _T_8672 = _T_8382 & _T_8380; // @[CLG.scala 26:31]
  assign _T_8673 = io_g[59]; // @[CLG.scala 18:18]
  assign _T_8674 = io_a[59]; // @[CLG.scala 19:18]
  assign _T_8967 = _T_8671 & _T_8674; // @[CLG.scala 26:21]
  assign _T_8968 = _T_8673 | _T_8967; // @[CLG.scala 26:11]
  assign _T_8969 = _T_8674 & _T_8672; // @[CLG.scala 26:31]
  assign _T_8970 = io_g[60]; // @[CLG.scala 18:18]
  assign _T_8971 = io_a[60]; // @[CLG.scala 19:18]
  assign _T_9269 = _T_8968 & _T_8971; // @[CLG.scala 26:21]
  assign _T_9270 = _T_8970 | _T_9269; // @[CLG.scala 26:11]
  assign _T_9271 = _T_8971 & _T_8969; // @[CLG.scala 26:31]
  assign _T_9272 = io_g[61]; // @[CLG.scala 18:18]
  assign _T_9273 = io_a[61]; // @[CLG.scala 19:18]
  assign _T_9576 = _T_9270 & _T_9273; // @[CLG.scala 26:21]
  assign _T_9577 = _T_9272 | _T_9576; // @[CLG.scala 26:11]
  assign _T_9578 = _T_9273 & _T_9271; // @[CLG.scala 26:31]
  assign _T_9579 = io_g[62]; // @[CLG.scala 18:18]
  assign _T_9580 = io_a[62]; // @[CLG.scala 19:18]
  assign _T_9888 = _T_9577 & _T_9580; // @[CLG.scala 26:21]
  assign _T_9889 = _T_9579 | _T_9888; // @[CLG.scala 26:11]
  assign _T_9890 = _T_9580 & _T_9578; // @[CLG.scala 26:31]
  assign _T_9891 = io_g[63]; // @[CLG.scala 18:18]
  assign _T_9892 = io_a[63]; // @[CLG.scala 19:18]
  assign _T_10205 = _T_9889 & _T_9892; // @[CLG.scala 26:21]
  assign _T_10206 = _T_9891 | _T_10205; // @[CLG.scala 26:11]
  assign _T_10207 = _T_9892 & _T_9890; // @[CLG.scala 26:31]
  assign _T_10208 = _T_1 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_0 = _T | _T_10208; // @[CLG.scala 41:12]
  assign _T_10209 = _T_8 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_1 = _T_7 | _T_10209; // @[CLG.scala 41:12]
  assign _T_10210 = _T_20 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_2 = _T_19 | _T_10210; // @[CLG.scala 41:12]
  assign _T_10211 = _T_37 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_3 = _T_36 | _T_10211; // @[CLG.scala 41:12]
  assign _T_10212 = _T_59 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_4 = _T_58 | _T_10212; // @[CLG.scala 41:12]
  assign _T_10213 = _T_86 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_5 = _T_85 | _T_10213; // @[CLG.scala 41:12]
  assign _T_10214 = _T_118 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_6 = _T_117 | _T_10214; // @[CLG.scala 41:12]
  assign _T_10215 = _T_155 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_7 = _T_154 | _T_10215; // @[CLG.scala 41:12]
  assign _T_10216 = _T_197 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_8 = _T_196 | _T_10216; // @[CLG.scala 41:12]
  assign _T_10217 = _T_244 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_9 = _T_243 | _T_10217; // @[CLG.scala 41:12]
  assign _T_10218 = _T_296 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_10 = _T_295 | _T_10218; // @[CLG.scala 41:12]
  assign _T_10219 = _T_353 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_11 = _T_352 | _T_10219; // @[CLG.scala 41:12]
  assign _T_10220 = _T_415 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_12 = _T_414 | _T_10220; // @[CLG.scala 41:12]
  assign _T_10221 = _T_482 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_13 = _T_481 | _T_10221; // @[CLG.scala 41:12]
  assign _T_10222 = _T_554 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_14 = _T_553 | _T_10222; // @[CLG.scala 41:12]
  assign _T_10223 = _T_631 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_15 = _T_630 | _T_10223; // @[CLG.scala 41:12]
  assign _T_10224 = _T_713 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_16 = _T_712 | _T_10224; // @[CLG.scala 41:12]
  assign _T_10225 = _T_800 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_17 = _T_799 | _T_10225; // @[CLG.scala 41:12]
  assign _T_10226 = _T_892 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_18 = _T_891 | _T_10226; // @[CLG.scala 41:12]
  assign _T_10227 = _T_989 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_19 = _T_988 | _T_10227; // @[CLG.scala 41:12]
  assign _T_10228 = _T_1091 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_20 = _T_1090 | _T_10228; // @[CLG.scala 41:12]
  assign _T_10229 = _T_1198 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_21 = _T_1197 | _T_10229; // @[CLG.scala 41:12]
  assign _T_10230 = _T_1310 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_22 = _T_1309 | _T_10230; // @[CLG.scala 41:12]
  assign _T_10231 = _T_1427 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_23 = _T_1426 | _T_10231; // @[CLG.scala 41:12]
  assign _T_10232 = _T_1549 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_24 = _T_1548 | _T_10232; // @[CLG.scala 41:12]
  assign _T_10233 = _T_1676 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_25 = _T_1675 | _T_10233; // @[CLG.scala 41:12]
  assign _T_10234 = _T_1808 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_26 = _T_1807 | _T_10234; // @[CLG.scala 41:12]
  assign _T_10235 = _T_1945 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_27 = _T_1944 | _T_10235; // @[CLG.scala 41:12]
  assign _T_10236 = _T_2087 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_28 = _T_2086 | _T_10236; // @[CLG.scala 41:12]
  assign _T_10237 = _T_2234 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_29 = _T_2233 | _T_10237; // @[CLG.scala 41:12]
  assign _T_10238 = _T_2386 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_30 = _T_2385 | _T_10238; // @[CLG.scala 41:12]
  assign _T_10239 = _T_2543 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_31 = _T_2542 | _T_10239; // @[CLG.scala 41:12]
  assign _T_10240 = _T_2705 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_32 = _T_2704 | _T_10240; // @[CLG.scala 41:12]
  assign _T_10241 = _T_2872 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_33 = _T_2871 | _T_10241; // @[CLG.scala 41:12]
  assign _T_10242 = _T_3044 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_34 = _T_3043 | _T_10242; // @[CLG.scala 41:12]
  assign _T_10243 = _T_3221 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_35 = _T_3220 | _T_10243; // @[CLG.scala 41:12]
  assign _T_10244 = _T_3403 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_36 = _T_3402 | _T_10244; // @[CLG.scala 41:12]
  assign _T_10245 = _T_3590 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_37 = _T_3589 | _T_10245; // @[CLG.scala 41:12]
  assign _T_10246 = _T_3782 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_38 = _T_3781 | _T_10246; // @[CLG.scala 41:12]
  assign _T_10247 = _T_3979 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_39 = _T_3978 | _T_10247; // @[CLG.scala 41:12]
  assign _T_10248 = _T_4181 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_40 = _T_4180 | _T_10248; // @[CLG.scala 41:12]
  assign _T_10249 = _T_4388 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_41 = _T_4387 | _T_10249; // @[CLG.scala 41:12]
  assign _T_10250 = _T_4600 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_42 = _T_4599 | _T_10250; // @[CLG.scala 41:12]
  assign _T_10251 = _T_4817 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_43 = _T_4816 | _T_10251; // @[CLG.scala 41:12]
  assign _T_10252 = _T_5039 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_44 = _T_5038 | _T_10252; // @[CLG.scala 41:12]
  assign _T_10253 = _T_5266 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_45 = _T_5265 | _T_10253; // @[CLG.scala 41:12]
  assign _T_10254 = _T_5498 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_46 = _T_5497 | _T_10254; // @[CLG.scala 41:12]
  assign _T_10255 = _T_5735 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_47 = _T_5734 | _T_10255; // @[CLG.scala 41:12]
  assign _T_10256 = _T_5977 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_48 = _T_5976 | _T_10256; // @[CLG.scala 41:12]
  assign _T_10257 = _T_6224 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_49 = _T_6223 | _T_10257; // @[CLG.scala 41:12]
  assign _T_10258 = _T_6476 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_50 = _T_6475 | _T_10258; // @[CLG.scala 41:12]
  assign _T_10259 = _T_6733 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_51 = _T_6732 | _T_10259; // @[CLG.scala 41:12]
  assign _T_10260 = _T_6995 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_52 = _T_6994 | _T_10260; // @[CLG.scala 41:12]
  assign _T_10261 = _T_7262 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_53 = _T_7261 | _T_10261; // @[CLG.scala 41:12]
  assign _T_10262 = _T_7534 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_54 = _T_7533 | _T_10262; // @[CLG.scala 41:12]
  assign _T_10263 = _T_7811 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_55 = _T_7810 | _T_10263; // @[CLG.scala 41:12]
  assign _T_10264 = _T_8093 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_56 = _T_8092 | _T_10264; // @[CLG.scala 41:12]
  assign _T_10265 = _T_8380 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_57 = _T_8379 | _T_10265; // @[CLG.scala 41:12]
  assign _T_10266 = _T_8672 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_58 = _T_8671 | _T_10266; // @[CLG.scala 41:12]
  assign _T_10267 = _T_8969 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_59 = _T_8968 | _T_10267; // @[CLG.scala 41:12]
  assign _T_10268 = _T_9271 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_60 = _T_9270 | _T_10268; // @[CLG.scala 41:12]
  assign _T_10269 = _T_9578 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_61 = _T_9577 | _T_10269; // @[CLG.scala 41:12]
  assign _T_10270 = _T_9890 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_62 = _T_9889 | _T_10270; // @[CLG.scala 41:12]
  assign _T_10271 = _T_10207 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_63 = _T_10206 | _T_10271; // @[CLG.scala 41:12]
  assign _T_10279 = {c_bit_7,c_bit_6,c_bit_5,c_bit_4,c_bit_3,c_bit_2,c_bit_1,c_bit_0}; // @[CLG.scala 43:32]
  assign _T_10287 = {c_bit_15,c_bit_14,c_bit_13,c_bit_12,c_bit_11,c_bit_10,c_bit_9,c_bit_8,_T_10279}; // @[CLG.scala 43:32]
  assign _T_10294 = {c_bit_23,c_bit_22,c_bit_21,c_bit_20,c_bit_19,c_bit_18,c_bit_17,c_bit_16}; // @[CLG.scala 43:32]
  assign _T_10303 = {c_bit_31,c_bit_30,c_bit_29,c_bit_28,c_bit_27,c_bit_26,c_bit_25,c_bit_24,_T_10294,_T_10287}; // @[CLG.scala 43:32]
  assign _T_10310 = {c_bit_39,c_bit_38,c_bit_37,c_bit_36,c_bit_35,c_bit_34,c_bit_33,c_bit_32}; // @[CLG.scala 43:32]
  assign _T_10318 = {c_bit_47,c_bit_46,c_bit_45,c_bit_44,c_bit_43,c_bit_42,c_bit_41,c_bit_40,_T_10310}; // @[CLG.scala 43:32]
  assign _T_10325 = {c_bit_55,c_bit_54,c_bit_53,c_bit_52,c_bit_51,c_bit_50,c_bit_49,c_bit_48}; // @[CLG.scala 43:32]
  assign _T_10334 = {c_bit_63,c_bit_62,c_bit_61,c_bit_60,c_bit_59,c_bit_58,c_bit_57,c_bit_56,_T_10325,_T_10318}; // @[CLG.scala 43:32]
  assign io_c = {_T_10334,_T_10303}; // @[CLG.scala 43:8]
  assign io_G = _T_9891 | _T_10205; // @[CLG.scala 46:8]
  assign io_A = _T_9892 & _T_9890; // @[CLG.scala 47:8]
endmodule
module CLA(
  input         clock,
  input         reset,
  input  [63:0] io_x,
  input  [63:0] io_y,
  input         io_cin,
  output [63:0] io_s,
  output        io_cout,
  output        io_G,
  output        io_A
);
  wire  GPA1_io_x; // @[CLA.scala 25:21]
  wire  GPA1_io_y; // @[CLA.scala 25:21]
  wire  GPA1_io_g; // @[CLA.scala 25:21]
  wire  GPA1_io_p; // @[CLA.scala 25:21]
  wire  GPA1_io_a; // @[CLA.scala 25:21]
  wire  GPA1_1_io_x; // @[CLA.scala 25:21]
  wire  GPA1_1_io_y; // @[CLA.scala 25:21]
  wire  GPA1_1_io_g; // @[CLA.scala 25:21]
  wire  GPA1_1_io_p; // @[CLA.scala 25:21]
  wire  GPA1_1_io_a; // @[CLA.scala 25:21]
  wire  GPA1_2_io_x; // @[CLA.scala 25:21]
  wire  GPA1_2_io_y; // @[CLA.scala 25:21]
  wire  GPA1_2_io_g; // @[CLA.scala 25:21]
  wire  GPA1_2_io_p; // @[CLA.scala 25:21]
  wire  GPA1_2_io_a; // @[CLA.scala 25:21]
  wire  GPA1_3_io_x; // @[CLA.scala 25:21]
  wire  GPA1_3_io_y; // @[CLA.scala 25:21]
  wire  GPA1_3_io_g; // @[CLA.scala 25:21]
  wire  GPA1_3_io_p; // @[CLA.scala 25:21]
  wire  GPA1_3_io_a; // @[CLA.scala 25:21]
  wire  GPA1_4_io_x; // @[CLA.scala 25:21]
  wire  GPA1_4_io_y; // @[CLA.scala 25:21]
  wire  GPA1_4_io_g; // @[CLA.scala 25:21]
  wire  GPA1_4_io_p; // @[CLA.scala 25:21]
  wire  GPA1_4_io_a; // @[CLA.scala 25:21]
  wire  GPA1_5_io_x; // @[CLA.scala 25:21]
  wire  GPA1_5_io_y; // @[CLA.scala 25:21]
  wire  GPA1_5_io_g; // @[CLA.scala 25:21]
  wire  GPA1_5_io_p; // @[CLA.scala 25:21]
  wire  GPA1_5_io_a; // @[CLA.scala 25:21]
  wire  GPA1_6_io_x; // @[CLA.scala 25:21]
  wire  GPA1_6_io_y; // @[CLA.scala 25:21]
  wire  GPA1_6_io_g; // @[CLA.scala 25:21]
  wire  GPA1_6_io_p; // @[CLA.scala 25:21]
  wire  GPA1_6_io_a; // @[CLA.scala 25:21]
  wire  GPA1_7_io_x; // @[CLA.scala 25:21]
  wire  GPA1_7_io_y; // @[CLA.scala 25:21]
  wire  GPA1_7_io_g; // @[CLA.scala 25:21]
  wire  GPA1_7_io_p; // @[CLA.scala 25:21]
  wire  GPA1_7_io_a; // @[CLA.scala 25:21]
  wire  GPA1_8_io_x; // @[CLA.scala 25:21]
  wire  GPA1_8_io_y; // @[CLA.scala 25:21]
  wire  GPA1_8_io_g; // @[CLA.scala 25:21]
  wire  GPA1_8_io_p; // @[CLA.scala 25:21]
  wire  GPA1_8_io_a; // @[CLA.scala 25:21]
  wire  GPA1_9_io_x; // @[CLA.scala 25:21]
  wire  GPA1_9_io_y; // @[CLA.scala 25:21]
  wire  GPA1_9_io_g; // @[CLA.scala 25:21]
  wire  GPA1_9_io_p; // @[CLA.scala 25:21]
  wire  GPA1_9_io_a; // @[CLA.scala 25:21]
  wire  GPA1_10_io_x; // @[CLA.scala 25:21]
  wire  GPA1_10_io_y; // @[CLA.scala 25:21]
  wire  GPA1_10_io_g; // @[CLA.scala 25:21]
  wire  GPA1_10_io_p; // @[CLA.scala 25:21]
  wire  GPA1_10_io_a; // @[CLA.scala 25:21]
  wire  GPA1_11_io_x; // @[CLA.scala 25:21]
  wire  GPA1_11_io_y; // @[CLA.scala 25:21]
  wire  GPA1_11_io_g; // @[CLA.scala 25:21]
  wire  GPA1_11_io_p; // @[CLA.scala 25:21]
  wire  GPA1_11_io_a; // @[CLA.scala 25:21]
  wire  GPA1_12_io_x; // @[CLA.scala 25:21]
  wire  GPA1_12_io_y; // @[CLA.scala 25:21]
  wire  GPA1_12_io_g; // @[CLA.scala 25:21]
  wire  GPA1_12_io_p; // @[CLA.scala 25:21]
  wire  GPA1_12_io_a; // @[CLA.scala 25:21]
  wire  GPA1_13_io_x; // @[CLA.scala 25:21]
  wire  GPA1_13_io_y; // @[CLA.scala 25:21]
  wire  GPA1_13_io_g; // @[CLA.scala 25:21]
  wire  GPA1_13_io_p; // @[CLA.scala 25:21]
  wire  GPA1_13_io_a; // @[CLA.scala 25:21]
  wire  GPA1_14_io_x; // @[CLA.scala 25:21]
  wire  GPA1_14_io_y; // @[CLA.scala 25:21]
  wire  GPA1_14_io_g; // @[CLA.scala 25:21]
  wire  GPA1_14_io_p; // @[CLA.scala 25:21]
  wire  GPA1_14_io_a; // @[CLA.scala 25:21]
  wire  GPA1_15_io_x; // @[CLA.scala 25:21]
  wire  GPA1_15_io_y; // @[CLA.scala 25:21]
  wire  GPA1_15_io_g; // @[CLA.scala 25:21]
  wire  GPA1_15_io_p; // @[CLA.scala 25:21]
  wire  GPA1_15_io_a; // @[CLA.scala 25:21]
  wire  GPA1_16_io_x; // @[CLA.scala 25:21]
  wire  GPA1_16_io_y; // @[CLA.scala 25:21]
  wire  GPA1_16_io_g; // @[CLA.scala 25:21]
  wire  GPA1_16_io_p; // @[CLA.scala 25:21]
  wire  GPA1_16_io_a; // @[CLA.scala 25:21]
  wire  GPA1_17_io_x; // @[CLA.scala 25:21]
  wire  GPA1_17_io_y; // @[CLA.scala 25:21]
  wire  GPA1_17_io_g; // @[CLA.scala 25:21]
  wire  GPA1_17_io_p; // @[CLA.scala 25:21]
  wire  GPA1_17_io_a; // @[CLA.scala 25:21]
  wire  GPA1_18_io_x; // @[CLA.scala 25:21]
  wire  GPA1_18_io_y; // @[CLA.scala 25:21]
  wire  GPA1_18_io_g; // @[CLA.scala 25:21]
  wire  GPA1_18_io_p; // @[CLA.scala 25:21]
  wire  GPA1_18_io_a; // @[CLA.scala 25:21]
  wire  GPA1_19_io_x; // @[CLA.scala 25:21]
  wire  GPA1_19_io_y; // @[CLA.scala 25:21]
  wire  GPA1_19_io_g; // @[CLA.scala 25:21]
  wire  GPA1_19_io_p; // @[CLA.scala 25:21]
  wire  GPA1_19_io_a; // @[CLA.scala 25:21]
  wire  GPA1_20_io_x; // @[CLA.scala 25:21]
  wire  GPA1_20_io_y; // @[CLA.scala 25:21]
  wire  GPA1_20_io_g; // @[CLA.scala 25:21]
  wire  GPA1_20_io_p; // @[CLA.scala 25:21]
  wire  GPA1_20_io_a; // @[CLA.scala 25:21]
  wire  GPA1_21_io_x; // @[CLA.scala 25:21]
  wire  GPA1_21_io_y; // @[CLA.scala 25:21]
  wire  GPA1_21_io_g; // @[CLA.scala 25:21]
  wire  GPA1_21_io_p; // @[CLA.scala 25:21]
  wire  GPA1_21_io_a; // @[CLA.scala 25:21]
  wire  GPA1_22_io_x; // @[CLA.scala 25:21]
  wire  GPA1_22_io_y; // @[CLA.scala 25:21]
  wire  GPA1_22_io_g; // @[CLA.scala 25:21]
  wire  GPA1_22_io_p; // @[CLA.scala 25:21]
  wire  GPA1_22_io_a; // @[CLA.scala 25:21]
  wire  GPA1_23_io_x; // @[CLA.scala 25:21]
  wire  GPA1_23_io_y; // @[CLA.scala 25:21]
  wire  GPA1_23_io_g; // @[CLA.scala 25:21]
  wire  GPA1_23_io_p; // @[CLA.scala 25:21]
  wire  GPA1_23_io_a; // @[CLA.scala 25:21]
  wire  GPA1_24_io_x; // @[CLA.scala 25:21]
  wire  GPA1_24_io_y; // @[CLA.scala 25:21]
  wire  GPA1_24_io_g; // @[CLA.scala 25:21]
  wire  GPA1_24_io_p; // @[CLA.scala 25:21]
  wire  GPA1_24_io_a; // @[CLA.scala 25:21]
  wire  GPA1_25_io_x; // @[CLA.scala 25:21]
  wire  GPA1_25_io_y; // @[CLA.scala 25:21]
  wire  GPA1_25_io_g; // @[CLA.scala 25:21]
  wire  GPA1_25_io_p; // @[CLA.scala 25:21]
  wire  GPA1_25_io_a; // @[CLA.scala 25:21]
  wire  GPA1_26_io_x; // @[CLA.scala 25:21]
  wire  GPA1_26_io_y; // @[CLA.scala 25:21]
  wire  GPA1_26_io_g; // @[CLA.scala 25:21]
  wire  GPA1_26_io_p; // @[CLA.scala 25:21]
  wire  GPA1_26_io_a; // @[CLA.scala 25:21]
  wire  GPA1_27_io_x; // @[CLA.scala 25:21]
  wire  GPA1_27_io_y; // @[CLA.scala 25:21]
  wire  GPA1_27_io_g; // @[CLA.scala 25:21]
  wire  GPA1_27_io_p; // @[CLA.scala 25:21]
  wire  GPA1_27_io_a; // @[CLA.scala 25:21]
  wire  GPA1_28_io_x; // @[CLA.scala 25:21]
  wire  GPA1_28_io_y; // @[CLA.scala 25:21]
  wire  GPA1_28_io_g; // @[CLA.scala 25:21]
  wire  GPA1_28_io_p; // @[CLA.scala 25:21]
  wire  GPA1_28_io_a; // @[CLA.scala 25:21]
  wire  GPA1_29_io_x; // @[CLA.scala 25:21]
  wire  GPA1_29_io_y; // @[CLA.scala 25:21]
  wire  GPA1_29_io_g; // @[CLA.scala 25:21]
  wire  GPA1_29_io_p; // @[CLA.scala 25:21]
  wire  GPA1_29_io_a; // @[CLA.scala 25:21]
  wire  GPA1_30_io_x; // @[CLA.scala 25:21]
  wire  GPA1_30_io_y; // @[CLA.scala 25:21]
  wire  GPA1_30_io_g; // @[CLA.scala 25:21]
  wire  GPA1_30_io_p; // @[CLA.scala 25:21]
  wire  GPA1_30_io_a; // @[CLA.scala 25:21]
  wire  GPA1_31_io_x; // @[CLA.scala 25:21]
  wire  GPA1_31_io_y; // @[CLA.scala 25:21]
  wire  GPA1_31_io_g; // @[CLA.scala 25:21]
  wire  GPA1_31_io_p; // @[CLA.scala 25:21]
  wire  GPA1_31_io_a; // @[CLA.scala 25:21]
  wire  GPA1_32_io_x; // @[CLA.scala 25:21]
  wire  GPA1_32_io_y; // @[CLA.scala 25:21]
  wire  GPA1_32_io_g; // @[CLA.scala 25:21]
  wire  GPA1_32_io_p; // @[CLA.scala 25:21]
  wire  GPA1_32_io_a; // @[CLA.scala 25:21]
  wire  GPA1_33_io_x; // @[CLA.scala 25:21]
  wire  GPA1_33_io_y; // @[CLA.scala 25:21]
  wire  GPA1_33_io_g; // @[CLA.scala 25:21]
  wire  GPA1_33_io_p; // @[CLA.scala 25:21]
  wire  GPA1_33_io_a; // @[CLA.scala 25:21]
  wire  GPA1_34_io_x; // @[CLA.scala 25:21]
  wire  GPA1_34_io_y; // @[CLA.scala 25:21]
  wire  GPA1_34_io_g; // @[CLA.scala 25:21]
  wire  GPA1_34_io_p; // @[CLA.scala 25:21]
  wire  GPA1_34_io_a; // @[CLA.scala 25:21]
  wire  GPA1_35_io_x; // @[CLA.scala 25:21]
  wire  GPA1_35_io_y; // @[CLA.scala 25:21]
  wire  GPA1_35_io_g; // @[CLA.scala 25:21]
  wire  GPA1_35_io_p; // @[CLA.scala 25:21]
  wire  GPA1_35_io_a; // @[CLA.scala 25:21]
  wire  GPA1_36_io_x; // @[CLA.scala 25:21]
  wire  GPA1_36_io_y; // @[CLA.scala 25:21]
  wire  GPA1_36_io_g; // @[CLA.scala 25:21]
  wire  GPA1_36_io_p; // @[CLA.scala 25:21]
  wire  GPA1_36_io_a; // @[CLA.scala 25:21]
  wire  GPA1_37_io_x; // @[CLA.scala 25:21]
  wire  GPA1_37_io_y; // @[CLA.scala 25:21]
  wire  GPA1_37_io_g; // @[CLA.scala 25:21]
  wire  GPA1_37_io_p; // @[CLA.scala 25:21]
  wire  GPA1_37_io_a; // @[CLA.scala 25:21]
  wire  GPA1_38_io_x; // @[CLA.scala 25:21]
  wire  GPA1_38_io_y; // @[CLA.scala 25:21]
  wire  GPA1_38_io_g; // @[CLA.scala 25:21]
  wire  GPA1_38_io_p; // @[CLA.scala 25:21]
  wire  GPA1_38_io_a; // @[CLA.scala 25:21]
  wire  GPA1_39_io_x; // @[CLA.scala 25:21]
  wire  GPA1_39_io_y; // @[CLA.scala 25:21]
  wire  GPA1_39_io_g; // @[CLA.scala 25:21]
  wire  GPA1_39_io_p; // @[CLA.scala 25:21]
  wire  GPA1_39_io_a; // @[CLA.scala 25:21]
  wire  GPA1_40_io_x; // @[CLA.scala 25:21]
  wire  GPA1_40_io_y; // @[CLA.scala 25:21]
  wire  GPA1_40_io_g; // @[CLA.scala 25:21]
  wire  GPA1_40_io_p; // @[CLA.scala 25:21]
  wire  GPA1_40_io_a; // @[CLA.scala 25:21]
  wire  GPA1_41_io_x; // @[CLA.scala 25:21]
  wire  GPA1_41_io_y; // @[CLA.scala 25:21]
  wire  GPA1_41_io_g; // @[CLA.scala 25:21]
  wire  GPA1_41_io_p; // @[CLA.scala 25:21]
  wire  GPA1_41_io_a; // @[CLA.scala 25:21]
  wire  GPA1_42_io_x; // @[CLA.scala 25:21]
  wire  GPA1_42_io_y; // @[CLA.scala 25:21]
  wire  GPA1_42_io_g; // @[CLA.scala 25:21]
  wire  GPA1_42_io_p; // @[CLA.scala 25:21]
  wire  GPA1_42_io_a; // @[CLA.scala 25:21]
  wire  GPA1_43_io_x; // @[CLA.scala 25:21]
  wire  GPA1_43_io_y; // @[CLA.scala 25:21]
  wire  GPA1_43_io_g; // @[CLA.scala 25:21]
  wire  GPA1_43_io_p; // @[CLA.scala 25:21]
  wire  GPA1_43_io_a; // @[CLA.scala 25:21]
  wire  GPA1_44_io_x; // @[CLA.scala 25:21]
  wire  GPA1_44_io_y; // @[CLA.scala 25:21]
  wire  GPA1_44_io_g; // @[CLA.scala 25:21]
  wire  GPA1_44_io_p; // @[CLA.scala 25:21]
  wire  GPA1_44_io_a; // @[CLA.scala 25:21]
  wire  GPA1_45_io_x; // @[CLA.scala 25:21]
  wire  GPA1_45_io_y; // @[CLA.scala 25:21]
  wire  GPA1_45_io_g; // @[CLA.scala 25:21]
  wire  GPA1_45_io_p; // @[CLA.scala 25:21]
  wire  GPA1_45_io_a; // @[CLA.scala 25:21]
  wire  GPA1_46_io_x; // @[CLA.scala 25:21]
  wire  GPA1_46_io_y; // @[CLA.scala 25:21]
  wire  GPA1_46_io_g; // @[CLA.scala 25:21]
  wire  GPA1_46_io_p; // @[CLA.scala 25:21]
  wire  GPA1_46_io_a; // @[CLA.scala 25:21]
  wire  GPA1_47_io_x; // @[CLA.scala 25:21]
  wire  GPA1_47_io_y; // @[CLA.scala 25:21]
  wire  GPA1_47_io_g; // @[CLA.scala 25:21]
  wire  GPA1_47_io_p; // @[CLA.scala 25:21]
  wire  GPA1_47_io_a; // @[CLA.scala 25:21]
  wire  GPA1_48_io_x; // @[CLA.scala 25:21]
  wire  GPA1_48_io_y; // @[CLA.scala 25:21]
  wire  GPA1_48_io_g; // @[CLA.scala 25:21]
  wire  GPA1_48_io_p; // @[CLA.scala 25:21]
  wire  GPA1_48_io_a; // @[CLA.scala 25:21]
  wire  GPA1_49_io_x; // @[CLA.scala 25:21]
  wire  GPA1_49_io_y; // @[CLA.scala 25:21]
  wire  GPA1_49_io_g; // @[CLA.scala 25:21]
  wire  GPA1_49_io_p; // @[CLA.scala 25:21]
  wire  GPA1_49_io_a; // @[CLA.scala 25:21]
  wire  GPA1_50_io_x; // @[CLA.scala 25:21]
  wire  GPA1_50_io_y; // @[CLA.scala 25:21]
  wire  GPA1_50_io_g; // @[CLA.scala 25:21]
  wire  GPA1_50_io_p; // @[CLA.scala 25:21]
  wire  GPA1_50_io_a; // @[CLA.scala 25:21]
  wire  GPA1_51_io_x; // @[CLA.scala 25:21]
  wire  GPA1_51_io_y; // @[CLA.scala 25:21]
  wire  GPA1_51_io_g; // @[CLA.scala 25:21]
  wire  GPA1_51_io_p; // @[CLA.scala 25:21]
  wire  GPA1_51_io_a; // @[CLA.scala 25:21]
  wire  GPA1_52_io_x; // @[CLA.scala 25:21]
  wire  GPA1_52_io_y; // @[CLA.scala 25:21]
  wire  GPA1_52_io_g; // @[CLA.scala 25:21]
  wire  GPA1_52_io_p; // @[CLA.scala 25:21]
  wire  GPA1_52_io_a; // @[CLA.scala 25:21]
  wire  GPA1_53_io_x; // @[CLA.scala 25:21]
  wire  GPA1_53_io_y; // @[CLA.scala 25:21]
  wire  GPA1_53_io_g; // @[CLA.scala 25:21]
  wire  GPA1_53_io_p; // @[CLA.scala 25:21]
  wire  GPA1_53_io_a; // @[CLA.scala 25:21]
  wire  GPA1_54_io_x; // @[CLA.scala 25:21]
  wire  GPA1_54_io_y; // @[CLA.scala 25:21]
  wire  GPA1_54_io_g; // @[CLA.scala 25:21]
  wire  GPA1_54_io_p; // @[CLA.scala 25:21]
  wire  GPA1_54_io_a; // @[CLA.scala 25:21]
  wire  GPA1_55_io_x; // @[CLA.scala 25:21]
  wire  GPA1_55_io_y; // @[CLA.scala 25:21]
  wire  GPA1_55_io_g; // @[CLA.scala 25:21]
  wire  GPA1_55_io_p; // @[CLA.scala 25:21]
  wire  GPA1_55_io_a; // @[CLA.scala 25:21]
  wire  GPA1_56_io_x; // @[CLA.scala 25:21]
  wire  GPA1_56_io_y; // @[CLA.scala 25:21]
  wire  GPA1_56_io_g; // @[CLA.scala 25:21]
  wire  GPA1_56_io_p; // @[CLA.scala 25:21]
  wire  GPA1_56_io_a; // @[CLA.scala 25:21]
  wire  GPA1_57_io_x; // @[CLA.scala 25:21]
  wire  GPA1_57_io_y; // @[CLA.scala 25:21]
  wire  GPA1_57_io_g; // @[CLA.scala 25:21]
  wire  GPA1_57_io_p; // @[CLA.scala 25:21]
  wire  GPA1_57_io_a; // @[CLA.scala 25:21]
  wire  GPA1_58_io_x; // @[CLA.scala 25:21]
  wire  GPA1_58_io_y; // @[CLA.scala 25:21]
  wire  GPA1_58_io_g; // @[CLA.scala 25:21]
  wire  GPA1_58_io_p; // @[CLA.scala 25:21]
  wire  GPA1_58_io_a; // @[CLA.scala 25:21]
  wire  GPA1_59_io_x; // @[CLA.scala 25:21]
  wire  GPA1_59_io_y; // @[CLA.scala 25:21]
  wire  GPA1_59_io_g; // @[CLA.scala 25:21]
  wire  GPA1_59_io_p; // @[CLA.scala 25:21]
  wire  GPA1_59_io_a; // @[CLA.scala 25:21]
  wire  GPA1_60_io_x; // @[CLA.scala 25:21]
  wire  GPA1_60_io_y; // @[CLA.scala 25:21]
  wire  GPA1_60_io_g; // @[CLA.scala 25:21]
  wire  GPA1_60_io_p; // @[CLA.scala 25:21]
  wire  GPA1_60_io_a; // @[CLA.scala 25:21]
  wire  GPA1_61_io_x; // @[CLA.scala 25:21]
  wire  GPA1_61_io_y; // @[CLA.scala 25:21]
  wire  GPA1_61_io_g; // @[CLA.scala 25:21]
  wire  GPA1_61_io_p; // @[CLA.scala 25:21]
  wire  GPA1_61_io_a; // @[CLA.scala 25:21]
  wire  GPA1_62_io_x; // @[CLA.scala 25:21]
  wire  GPA1_62_io_y; // @[CLA.scala 25:21]
  wire  GPA1_62_io_g; // @[CLA.scala 25:21]
  wire  GPA1_62_io_p; // @[CLA.scala 25:21]
  wire  GPA1_62_io_a; // @[CLA.scala 25:21]
  wire  GPA1_63_io_x; // @[CLA.scala 25:21]
  wire  GPA1_63_io_y; // @[CLA.scala 25:21]
  wire  GPA1_63_io_g; // @[CLA.scala 25:21]
  wire  GPA1_63_io_p; // @[CLA.scala 25:21]
  wire  GPA1_63_io_a; // @[CLA.scala 25:21]
  wire [63:0] CLG_io_g; // @[CLA.scala 32:19]
  wire [63:0] CLG_io_a; // @[CLA.scala 32:19]
  wire  CLG_io_cin; // @[CLA.scala 32:19]
  wire [63:0] CLG_io_c; // @[CLA.scala 32:19]
  wire  CLG_io_G; // @[CLA.scala 32:19]
  wire  CLG_io_A; // @[CLA.scala 32:19]
  wire  _T_128_1; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_0; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_3; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_2; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_5; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_4; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_7; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_6; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_135; // @[CLA.scala 33:46]
  wire  _T_128_9; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_8; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_11; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_10; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_13; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_12; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_15; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_14; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [15:0] _T_143; // @[CLA.scala 33:46]
  wire  _T_128_17; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_16; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_19; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_18; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_21; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_20; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_23; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_22; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_150; // @[CLA.scala 33:46]
  wire  _T_128_25; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_24; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_27; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_26; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_29; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_28; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_31; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_30; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [31:0] _T_159; // @[CLA.scala 33:46]
  wire  _T_128_33; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_32; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_35; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_34; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_37; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_36; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_39; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_38; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_166; // @[CLA.scala 33:46]
  wire  _T_128_41; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_40; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_43; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_42; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_45; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_44; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_47; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_46; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [15:0] _T_174; // @[CLA.scala 33:46]
  wire  _T_128_49; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_48; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_51; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_50; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_53; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_52; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_55; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_54; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_181; // @[CLA.scala 33:46]
  wire  _T_128_57; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_56; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_59; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_58; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_61; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_60; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_63; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_128_62; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [31:0] _T_190; // @[CLA.scala 33:46]
  wire  _T_192_1; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_0; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_3; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_2; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_5; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_4; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_7; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_6; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_199; // @[CLA.scala 34:46]
  wire  _T_192_9; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_8; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_11; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_10; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_13; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_12; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_15; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_14; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [15:0] _T_207; // @[CLA.scala 34:46]
  wire  _T_192_17; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_16; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_19; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_18; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_21; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_20; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_23; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_22; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_214; // @[CLA.scala 34:46]
  wire  _T_192_25; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_24; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_27; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_26; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_29; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_28; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_31; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_30; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [31:0] _T_223; // @[CLA.scala 34:46]
  wire  _T_192_33; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_32; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_35; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_34; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_37; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_36; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_39; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_38; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_230; // @[CLA.scala 34:46]
  wire  _T_192_41; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_40; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_43; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_42; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_45; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_44; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_47; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_46; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [15:0] _T_238; // @[CLA.scala 34:46]
  wire  _T_192_49; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_48; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_51; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_50; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_53; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_52; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_55; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_54; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_245; // @[CLA.scala 34:46]
  wire  _T_192_57; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_56; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_59; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_58; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_61; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_60; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_63; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_192_62; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [31:0] _T_254; // @[CLA.scala 34:46]
  wire  s_bit_0; // @[CLA.scala 41:14]
  wire  _T_256; // @[CLA.scala 43:12]
  wire  s_bit_1; // @[CLA.scala 43:22]
  wire  _T_257; // @[CLA.scala 43:12]
  wire  s_bit_2; // @[CLA.scala 43:22]
  wire  _T_258; // @[CLA.scala 43:12]
  wire  s_bit_3; // @[CLA.scala 43:22]
  wire  _T_259; // @[CLA.scala 43:12]
  wire  s_bit_4; // @[CLA.scala 43:22]
  wire  _T_260; // @[CLA.scala 43:12]
  wire  s_bit_5; // @[CLA.scala 43:22]
  wire  _T_261; // @[CLA.scala 43:12]
  wire  s_bit_6; // @[CLA.scala 43:22]
  wire  _T_262; // @[CLA.scala 43:12]
  wire  s_bit_7; // @[CLA.scala 43:22]
  wire  _T_263; // @[CLA.scala 43:12]
  wire  s_bit_8; // @[CLA.scala 43:22]
  wire  _T_264; // @[CLA.scala 43:12]
  wire  s_bit_9; // @[CLA.scala 43:22]
  wire  _T_265; // @[CLA.scala 43:12]
  wire  s_bit_10; // @[CLA.scala 43:22]
  wire  _T_266; // @[CLA.scala 43:12]
  wire  s_bit_11; // @[CLA.scala 43:22]
  wire  _T_267; // @[CLA.scala 43:12]
  wire  s_bit_12; // @[CLA.scala 43:22]
  wire  _T_268; // @[CLA.scala 43:12]
  wire  s_bit_13; // @[CLA.scala 43:22]
  wire  _T_269; // @[CLA.scala 43:12]
  wire  s_bit_14; // @[CLA.scala 43:22]
  wire  _T_270; // @[CLA.scala 43:12]
  wire  s_bit_15; // @[CLA.scala 43:22]
  wire  _T_271; // @[CLA.scala 43:12]
  wire  s_bit_16; // @[CLA.scala 43:22]
  wire  _T_272; // @[CLA.scala 43:12]
  wire  s_bit_17; // @[CLA.scala 43:22]
  wire  _T_273; // @[CLA.scala 43:12]
  wire  s_bit_18; // @[CLA.scala 43:22]
  wire  _T_274; // @[CLA.scala 43:12]
  wire  s_bit_19; // @[CLA.scala 43:22]
  wire  _T_275; // @[CLA.scala 43:12]
  wire  s_bit_20; // @[CLA.scala 43:22]
  wire  _T_276; // @[CLA.scala 43:12]
  wire  s_bit_21; // @[CLA.scala 43:22]
  wire  _T_277; // @[CLA.scala 43:12]
  wire  s_bit_22; // @[CLA.scala 43:22]
  wire  _T_278; // @[CLA.scala 43:12]
  wire  s_bit_23; // @[CLA.scala 43:22]
  wire  _T_279; // @[CLA.scala 43:12]
  wire  s_bit_24; // @[CLA.scala 43:22]
  wire  _T_280; // @[CLA.scala 43:12]
  wire  s_bit_25; // @[CLA.scala 43:22]
  wire  _T_281; // @[CLA.scala 43:12]
  wire  s_bit_26; // @[CLA.scala 43:22]
  wire  _T_282; // @[CLA.scala 43:12]
  wire  s_bit_27; // @[CLA.scala 43:22]
  wire  _T_283; // @[CLA.scala 43:12]
  wire  s_bit_28; // @[CLA.scala 43:22]
  wire  _T_284; // @[CLA.scala 43:12]
  wire  s_bit_29; // @[CLA.scala 43:22]
  wire  _T_285; // @[CLA.scala 43:12]
  wire  s_bit_30; // @[CLA.scala 43:22]
  wire  _T_286; // @[CLA.scala 43:12]
  wire  s_bit_31; // @[CLA.scala 43:22]
  wire  _T_287; // @[CLA.scala 43:12]
  wire  s_bit_32; // @[CLA.scala 43:22]
  wire  _T_288; // @[CLA.scala 43:12]
  wire  s_bit_33; // @[CLA.scala 43:22]
  wire  _T_289; // @[CLA.scala 43:12]
  wire  s_bit_34; // @[CLA.scala 43:22]
  wire  _T_290; // @[CLA.scala 43:12]
  wire  s_bit_35; // @[CLA.scala 43:22]
  wire  _T_291; // @[CLA.scala 43:12]
  wire  s_bit_36; // @[CLA.scala 43:22]
  wire  _T_292; // @[CLA.scala 43:12]
  wire  s_bit_37; // @[CLA.scala 43:22]
  wire  _T_293; // @[CLA.scala 43:12]
  wire  s_bit_38; // @[CLA.scala 43:22]
  wire  _T_294; // @[CLA.scala 43:12]
  wire  s_bit_39; // @[CLA.scala 43:22]
  wire  _T_295; // @[CLA.scala 43:12]
  wire  s_bit_40; // @[CLA.scala 43:22]
  wire  _T_296; // @[CLA.scala 43:12]
  wire  s_bit_41; // @[CLA.scala 43:22]
  wire  _T_297; // @[CLA.scala 43:12]
  wire  s_bit_42; // @[CLA.scala 43:22]
  wire  _T_298; // @[CLA.scala 43:12]
  wire  s_bit_43; // @[CLA.scala 43:22]
  wire  _T_299; // @[CLA.scala 43:12]
  wire  s_bit_44; // @[CLA.scala 43:22]
  wire  _T_300; // @[CLA.scala 43:12]
  wire  s_bit_45; // @[CLA.scala 43:22]
  wire  _T_301; // @[CLA.scala 43:12]
  wire  s_bit_46; // @[CLA.scala 43:22]
  wire  _T_302; // @[CLA.scala 43:12]
  wire  s_bit_47; // @[CLA.scala 43:22]
  wire  _T_303; // @[CLA.scala 43:12]
  wire  s_bit_48; // @[CLA.scala 43:22]
  wire  _T_304; // @[CLA.scala 43:12]
  wire  s_bit_49; // @[CLA.scala 43:22]
  wire  _T_305; // @[CLA.scala 43:12]
  wire  s_bit_50; // @[CLA.scala 43:22]
  wire  _T_306; // @[CLA.scala 43:12]
  wire  s_bit_51; // @[CLA.scala 43:22]
  wire  _T_307; // @[CLA.scala 43:12]
  wire  s_bit_52; // @[CLA.scala 43:22]
  wire  _T_308; // @[CLA.scala 43:12]
  wire  s_bit_53; // @[CLA.scala 43:22]
  wire  _T_309; // @[CLA.scala 43:12]
  wire  s_bit_54; // @[CLA.scala 43:22]
  wire  _T_310; // @[CLA.scala 43:12]
  wire  s_bit_55; // @[CLA.scala 43:22]
  wire  _T_311; // @[CLA.scala 43:12]
  wire  s_bit_56; // @[CLA.scala 43:22]
  wire  _T_312; // @[CLA.scala 43:12]
  wire  s_bit_57; // @[CLA.scala 43:22]
  wire  _T_313; // @[CLA.scala 43:12]
  wire  s_bit_58; // @[CLA.scala 43:22]
  wire  _T_314; // @[CLA.scala 43:12]
  wire  s_bit_59; // @[CLA.scala 43:22]
  wire  _T_315; // @[CLA.scala 43:12]
  wire  s_bit_60; // @[CLA.scala 43:22]
  wire  _T_316; // @[CLA.scala 43:12]
  wire  s_bit_61; // @[CLA.scala 43:22]
  wire  _T_317; // @[CLA.scala 43:12]
  wire  s_bit_62; // @[CLA.scala 43:22]
  wire  _T_318; // @[CLA.scala 43:12]
  wire  s_bit_63; // @[CLA.scala 43:22]
  wire [7:0] _T_326; // @[CLA.scala 46:32]
  wire [15:0] _T_334; // @[CLA.scala 46:32]
  wire [7:0] _T_341; // @[CLA.scala 46:32]
  wire [31:0] _T_350; // @[CLA.scala 46:32]
  wire [7:0] _T_357; // @[CLA.scala 46:32]
  wire [15:0] _T_365; // @[CLA.scala 46:32]
  wire [7:0] _T_372; // @[CLA.scala 46:32]
  wire [31:0] _T_381; // @[CLA.scala 46:32]
  GPA1 GPA1 ( // @[CLA.scala 25:21]
    .io_x(GPA1_io_x),
    .io_y(GPA1_io_y),
    .io_g(GPA1_io_g),
    .io_p(GPA1_io_p),
    .io_a(GPA1_io_a)
  );
  GPA1 GPA1_1 ( // @[CLA.scala 25:21]
    .io_x(GPA1_1_io_x),
    .io_y(GPA1_1_io_y),
    .io_g(GPA1_1_io_g),
    .io_p(GPA1_1_io_p),
    .io_a(GPA1_1_io_a)
  );
  GPA1 GPA1_2 ( // @[CLA.scala 25:21]
    .io_x(GPA1_2_io_x),
    .io_y(GPA1_2_io_y),
    .io_g(GPA1_2_io_g),
    .io_p(GPA1_2_io_p),
    .io_a(GPA1_2_io_a)
  );
  GPA1 GPA1_3 ( // @[CLA.scala 25:21]
    .io_x(GPA1_3_io_x),
    .io_y(GPA1_3_io_y),
    .io_g(GPA1_3_io_g),
    .io_p(GPA1_3_io_p),
    .io_a(GPA1_3_io_a)
  );
  GPA1 GPA1_4 ( // @[CLA.scala 25:21]
    .io_x(GPA1_4_io_x),
    .io_y(GPA1_4_io_y),
    .io_g(GPA1_4_io_g),
    .io_p(GPA1_4_io_p),
    .io_a(GPA1_4_io_a)
  );
  GPA1 GPA1_5 ( // @[CLA.scala 25:21]
    .io_x(GPA1_5_io_x),
    .io_y(GPA1_5_io_y),
    .io_g(GPA1_5_io_g),
    .io_p(GPA1_5_io_p),
    .io_a(GPA1_5_io_a)
  );
  GPA1 GPA1_6 ( // @[CLA.scala 25:21]
    .io_x(GPA1_6_io_x),
    .io_y(GPA1_6_io_y),
    .io_g(GPA1_6_io_g),
    .io_p(GPA1_6_io_p),
    .io_a(GPA1_6_io_a)
  );
  GPA1 GPA1_7 ( // @[CLA.scala 25:21]
    .io_x(GPA1_7_io_x),
    .io_y(GPA1_7_io_y),
    .io_g(GPA1_7_io_g),
    .io_p(GPA1_7_io_p),
    .io_a(GPA1_7_io_a)
  );
  GPA1 GPA1_8 ( // @[CLA.scala 25:21]
    .io_x(GPA1_8_io_x),
    .io_y(GPA1_8_io_y),
    .io_g(GPA1_8_io_g),
    .io_p(GPA1_8_io_p),
    .io_a(GPA1_8_io_a)
  );
  GPA1 GPA1_9 ( // @[CLA.scala 25:21]
    .io_x(GPA1_9_io_x),
    .io_y(GPA1_9_io_y),
    .io_g(GPA1_9_io_g),
    .io_p(GPA1_9_io_p),
    .io_a(GPA1_9_io_a)
  );
  GPA1 GPA1_10 ( // @[CLA.scala 25:21]
    .io_x(GPA1_10_io_x),
    .io_y(GPA1_10_io_y),
    .io_g(GPA1_10_io_g),
    .io_p(GPA1_10_io_p),
    .io_a(GPA1_10_io_a)
  );
  GPA1 GPA1_11 ( // @[CLA.scala 25:21]
    .io_x(GPA1_11_io_x),
    .io_y(GPA1_11_io_y),
    .io_g(GPA1_11_io_g),
    .io_p(GPA1_11_io_p),
    .io_a(GPA1_11_io_a)
  );
  GPA1 GPA1_12 ( // @[CLA.scala 25:21]
    .io_x(GPA1_12_io_x),
    .io_y(GPA1_12_io_y),
    .io_g(GPA1_12_io_g),
    .io_p(GPA1_12_io_p),
    .io_a(GPA1_12_io_a)
  );
  GPA1 GPA1_13 ( // @[CLA.scala 25:21]
    .io_x(GPA1_13_io_x),
    .io_y(GPA1_13_io_y),
    .io_g(GPA1_13_io_g),
    .io_p(GPA1_13_io_p),
    .io_a(GPA1_13_io_a)
  );
  GPA1 GPA1_14 ( // @[CLA.scala 25:21]
    .io_x(GPA1_14_io_x),
    .io_y(GPA1_14_io_y),
    .io_g(GPA1_14_io_g),
    .io_p(GPA1_14_io_p),
    .io_a(GPA1_14_io_a)
  );
  GPA1 GPA1_15 ( // @[CLA.scala 25:21]
    .io_x(GPA1_15_io_x),
    .io_y(GPA1_15_io_y),
    .io_g(GPA1_15_io_g),
    .io_p(GPA1_15_io_p),
    .io_a(GPA1_15_io_a)
  );
  GPA1 GPA1_16 ( // @[CLA.scala 25:21]
    .io_x(GPA1_16_io_x),
    .io_y(GPA1_16_io_y),
    .io_g(GPA1_16_io_g),
    .io_p(GPA1_16_io_p),
    .io_a(GPA1_16_io_a)
  );
  GPA1 GPA1_17 ( // @[CLA.scala 25:21]
    .io_x(GPA1_17_io_x),
    .io_y(GPA1_17_io_y),
    .io_g(GPA1_17_io_g),
    .io_p(GPA1_17_io_p),
    .io_a(GPA1_17_io_a)
  );
  GPA1 GPA1_18 ( // @[CLA.scala 25:21]
    .io_x(GPA1_18_io_x),
    .io_y(GPA1_18_io_y),
    .io_g(GPA1_18_io_g),
    .io_p(GPA1_18_io_p),
    .io_a(GPA1_18_io_a)
  );
  GPA1 GPA1_19 ( // @[CLA.scala 25:21]
    .io_x(GPA1_19_io_x),
    .io_y(GPA1_19_io_y),
    .io_g(GPA1_19_io_g),
    .io_p(GPA1_19_io_p),
    .io_a(GPA1_19_io_a)
  );
  GPA1 GPA1_20 ( // @[CLA.scala 25:21]
    .io_x(GPA1_20_io_x),
    .io_y(GPA1_20_io_y),
    .io_g(GPA1_20_io_g),
    .io_p(GPA1_20_io_p),
    .io_a(GPA1_20_io_a)
  );
  GPA1 GPA1_21 ( // @[CLA.scala 25:21]
    .io_x(GPA1_21_io_x),
    .io_y(GPA1_21_io_y),
    .io_g(GPA1_21_io_g),
    .io_p(GPA1_21_io_p),
    .io_a(GPA1_21_io_a)
  );
  GPA1 GPA1_22 ( // @[CLA.scala 25:21]
    .io_x(GPA1_22_io_x),
    .io_y(GPA1_22_io_y),
    .io_g(GPA1_22_io_g),
    .io_p(GPA1_22_io_p),
    .io_a(GPA1_22_io_a)
  );
  GPA1 GPA1_23 ( // @[CLA.scala 25:21]
    .io_x(GPA1_23_io_x),
    .io_y(GPA1_23_io_y),
    .io_g(GPA1_23_io_g),
    .io_p(GPA1_23_io_p),
    .io_a(GPA1_23_io_a)
  );
  GPA1 GPA1_24 ( // @[CLA.scala 25:21]
    .io_x(GPA1_24_io_x),
    .io_y(GPA1_24_io_y),
    .io_g(GPA1_24_io_g),
    .io_p(GPA1_24_io_p),
    .io_a(GPA1_24_io_a)
  );
  GPA1 GPA1_25 ( // @[CLA.scala 25:21]
    .io_x(GPA1_25_io_x),
    .io_y(GPA1_25_io_y),
    .io_g(GPA1_25_io_g),
    .io_p(GPA1_25_io_p),
    .io_a(GPA1_25_io_a)
  );
  GPA1 GPA1_26 ( // @[CLA.scala 25:21]
    .io_x(GPA1_26_io_x),
    .io_y(GPA1_26_io_y),
    .io_g(GPA1_26_io_g),
    .io_p(GPA1_26_io_p),
    .io_a(GPA1_26_io_a)
  );
  GPA1 GPA1_27 ( // @[CLA.scala 25:21]
    .io_x(GPA1_27_io_x),
    .io_y(GPA1_27_io_y),
    .io_g(GPA1_27_io_g),
    .io_p(GPA1_27_io_p),
    .io_a(GPA1_27_io_a)
  );
  GPA1 GPA1_28 ( // @[CLA.scala 25:21]
    .io_x(GPA1_28_io_x),
    .io_y(GPA1_28_io_y),
    .io_g(GPA1_28_io_g),
    .io_p(GPA1_28_io_p),
    .io_a(GPA1_28_io_a)
  );
  GPA1 GPA1_29 ( // @[CLA.scala 25:21]
    .io_x(GPA1_29_io_x),
    .io_y(GPA1_29_io_y),
    .io_g(GPA1_29_io_g),
    .io_p(GPA1_29_io_p),
    .io_a(GPA1_29_io_a)
  );
  GPA1 GPA1_30 ( // @[CLA.scala 25:21]
    .io_x(GPA1_30_io_x),
    .io_y(GPA1_30_io_y),
    .io_g(GPA1_30_io_g),
    .io_p(GPA1_30_io_p),
    .io_a(GPA1_30_io_a)
  );
  GPA1 GPA1_31 ( // @[CLA.scala 25:21]
    .io_x(GPA1_31_io_x),
    .io_y(GPA1_31_io_y),
    .io_g(GPA1_31_io_g),
    .io_p(GPA1_31_io_p),
    .io_a(GPA1_31_io_a)
  );
  GPA1 GPA1_32 ( // @[CLA.scala 25:21]
    .io_x(GPA1_32_io_x),
    .io_y(GPA1_32_io_y),
    .io_g(GPA1_32_io_g),
    .io_p(GPA1_32_io_p),
    .io_a(GPA1_32_io_a)
  );
  GPA1 GPA1_33 ( // @[CLA.scala 25:21]
    .io_x(GPA1_33_io_x),
    .io_y(GPA1_33_io_y),
    .io_g(GPA1_33_io_g),
    .io_p(GPA1_33_io_p),
    .io_a(GPA1_33_io_a)
  );
  GPA1 GPA1_34 ( // @[CLA.scala 25:21]
    .io_x(GPA1_34_io_x),
    .io_y(GPA1_34_io_y),
    .io_g(GPA1_34_io_g),
    .io_p(GPA1_34_io_p),
    .io_a(GPA1_34_io_a)
  );
  GPA1 GPA1_35 ( // @[CLA.scala 25:21]
    .io_x(GPA1_35_io_x),
    .io_y(GPA1_35_io_y),
    .io_g(GPA1_35_io_g),
    .io_p(GPA1_35_io_p),
    .io_a(GPA1_35_io_a)
  );
  GPA1 GPA1_36 ( // @[CLA.scala 25:21]
    .io_x(GPA1_36_io_x),
    .io_y(GPA1_36_io_y),
    .io_g(GPA1_36_io_g),
    .io_p(GPA1_36_io_p),
    .io_a(GPA1_36_io_a)
  );
  GPA1 GPA1_37 ( // @[CLA.scala 25:21]
    .io_x(GPA1_37_io_x),
    .io_y(GPA1_37_io_y),
    .io_g(GPA1_37_io_g),
    .io_p(GPA1_37_io_p),
    .io_a(GPA1_37_io_a)
  );
  GPA1 GPA1_38 ( // @[CLA.scala 25:21]
    .io_x(GPA1_38_io_x),
    .io_y(GPA1_38_io_y),
    .io_g(GPA1_38_io_g),
    .io_p(GPA1_38_io_p),
    .io_a(GPA1_38_io_a)
  );
  GPA1 GPA1_39 ( // @[CLA.scala 25:21]
    .io_x(GPA1_39_io_x),
    .io_y(GPA1_39_io_y),
    .io_g(GPA1_39_io_g),
    .io_p(GPA1_39_io_p),
    .io_a(GPA1_39_io_a)
  );
  GPA1 GPA1_40 ( // @[CLA.scala 25:21]
    .io_x(GPA1_40_io_x),
    .io_y(GPA1_40_io_y),
    .io_g(GPA1_40_io_g),
    .io_p(GPA1_40_io_p),
    .io_a(GPA1_40_io_a)
  );
  GPA1 GPA1_41 ( // @[CLA.scala 25:21]
    .io_x(GPA1_41_io_x),
    .io_y(GPA1_41_io_y),
    .io_g(GPA1_41_io_g),
    .io_p(GPA1_41_io_p),
    .io_a(GPA1_41_io_a)
  );
  GPA1 GPA1_42 ( // @[CLA.scala 25:21]
    .io_x(GPA1_42_io_x),
    .io_y(GPA1_42_io_y),
    .io_g(GPA1_42_io_g),
    .io_p(GPA1_42_io_p),
    .io_a(GPA1_42_io_a)
  );
  GPA1 GPA1_43 ( // @[CLA.scala 25:21]
    .io_x(GPA1_43_io_x),
    .io_y(GPA1_43_io_y),
    .io_g(GPA1_43_io_g),
    .io_p(GPA1_43_io_p),
    .io_a(GPA1_43_io_a)
  );
  GPA1 GPA1_44 ( // @[CLA.scala 25:21]
    .io_x(GPA1_44_io_x),
    .io_y(GPA1_44_io_y),
    .io_g(GPA1_44_io_g),
    .io_p(GPA1_44_io_p),
    .io_a(GPA1_44_io_a)
  );
  GPA1 GPA1_45 ( // @[CLA.scala 25:21]
    .io_x(GPA1_45_io_x),
    .io_y(GPA1_45_io_y),
    .io_g(GPA1_45_io_g),
    .io_p(GPA1_45_io_p),
    .io_a(GPA1_45_io_a)
  );
  GPA1 GPA1_46 ( // @[CLA.scala 25:21]
    .io_x(GPA1_46_io_x),
    .io_y(GPA1_46_io_y),
    .io_g(GPA1_46_io_g),
    .io_p(GPA1_46_io_p),
    .io_a(GPA1_46_io_a)
  );
  GPA1 GPA1_47 ( // @[CLA.scala 25:21]
    .io_x(GPA1_47_io_x),
    .io_y(GPA1_47_io_y),
    .io_g(GPA1_47_io_g),
    .io_p(GPA1_47_io_p),
    .io_a(GPA1_47_io_a)
  );
  GPA1 GPA1_48 ( // @[CLA.scala 25:21]
    .io_x(GPA1_48_io_x),
    .io_y(GPA1_48_io_y),
    .io_g(GPA1_48_io_g),
    .io_p(GPA1_48_io_p),
    .io_a(GPA1_48_io_a)
  );
  GPA1 GPA1_49 ( // @[CLA.scala 25:21]
    .io_x(GPA1_49_io_x),
    .io_y(GPA1_49_io_y),
    .io_g(GPA1_49_io_g),
    .io_p(GPA1_49_io_p),
    .io_a(GPA1_49_io_a)
  );
  GPA1 GPA1_50 ( // @[CLA.scala 25:21]
    .io_x(GPA1_50_io_x),
    .io_y(GPA1_50_io_y),
    .io_g(GPA1_50_io_g),
    .io_p(GPA1_50_io_p),
    .io_a(GPA1_50_io_a)
  );
  GPA1 GPA1_51 ( // @[CLA.scala 25:21]
    .io_x(GPA1_51_io_x),
    .io_y(GPA1_51_io_y),
    .io_g(GPA1_51_io_g),
    .io_p(GPA1_51_io_p),
    .io_a(GPA1_51_io_a)
  );
  GPA1 GPA1_52 ( // @[CLA.scala 25:21]
    .io_x(GPA1_52_io_x),
    .io_y(GPA1_52_io_y),
    .io_g(GPA1_52_io_g),
    .io_p(GPA1_52_io_p),
    .io_a(GPA1_52_io_a)
  );
  GPA1 GPA1_53 ( // @[CLA.scala 25:21]
    .io_x(GPA1_53_io_x),
    .io_y(GPA1_53_io_y),
    .io_g(GPA1_53_io_g),
    .io_p(GPA1_53_io_p),
    .io_a(GPA1_53_io_a)
  );
  GPA1 GPA1_54 ( // @[CLA.scala 25:21]
    .io_x(GPA1_54_io_x),
    .io_y(GPA1_54_io_y),
    .io_g(GPA1_54_io_g),
    .io_p(GPA1_54_io_p),
    .io_a(GPA1_54_io_a)
  );
  GPA1 GPA1_55 ( // @[CLA.scala 25:21]
    .io_x(GPA1_55_io_x),
    .io_y(GPA1_55_io_y),
    .io_g(GPA1_55_io_g),
    .io_p(GPA1_55_io_p),
    .io_a(GPA1_55_io_a)
  );
  GPA1 GPA1_56 ( // @[CLA.scala 25:21]
    .io_x(GPA1_56_io_x),
    .io_y(GPA1_56_io_y),
    .io_g(GPA1_56_io_g),
    .io_p(GPA1_56_io_p),
    .io_a(GPA1_56_io_a)
  );
  GPA1 GPA1_57 ( // @[CLA.scala 25:21]
    .io_x(GPA1_57_io_x),
    .io_y(GPA1_57_io_y),
    .io_g(GPA1_57_io_g),
    .io_p(GPA1_57_io_p),
    .io_a(GPA1_57_io_a)
  );
  GPA1 GPA1_58 ( // @[CLA.scala 25:21]
    .io_x(GPA1_58_io_x),
    .io_y(GPA1_58_io_y),
    .io_g(GPA1_58_io_g),
    .io_p(GPA1_58_io_p),
    .io_a(GPA1_58_io_a)
  );
  GPA1 GPA1_59 ( // @[CLA.scala 25:21]
    .io_x(GPA1_59_io_x),
    .io_y(GPA1_59_io_y),
    .io_g(GPA1_59_io_g),
    .io_p(GPA1_59_io_p),
    .io_a(GPA1_59_io_a)
  );
  GPA1 GPA1_60 ( // @[CLA.scala 25:21]
    .io_x(GPA1_60_io_x),
    .io_y(GPA1_60_io_y),
    .io_g(GPA1_60_io_g),
    .io_p(GPA1_60_io_p),
    .io_a(GPA1_60_io_a)
  );
  GPA1 GPA1_61 ( // @[CLA.scala 25:21]
    .io_x(GPA1_61_io_x),
    .io_y(GPA1_61_io_y),
    .io_g(GPA1_61_io_g),
    .io_p(GPA1_61_io_p),
    .io_a(GPA1_61_io_a)
  );
  GPA1 GPA1_62 ( // @[CLA.scala 25:21]
    .io_x(GPA1_62_io_x),
    .io_y(GPA1_62_io_y),
    .io_g(GPA1_62_io_g),
    .io_p(GPA1_62_io_p),
    .io_a(GPA1_62_io_a)
  );
  GPA1 GPA1_63 ( // @[CLA.scala 25:21]
    .io_x(GPA1_63_io_x),
    .io_y(GPA1_63_io_y),
    .io_g(GPA1_63_io_g),
    .io_p(GPA1_63_io_p),
    .io_a(GPA1_63_io_a)
  );
  CLG CLG ( // @[CLA.scala 32:19]
    .io_g(CLG_io_g),
    .io_a(CLG_io_a),
    .io_cin(CLG_io_cin),
    .io_c(CLG_io_c),
    .io_G(CLG_io_G),
    .io_A(CLG_io_A)
  );
  assign _T_128_1 = GPA1_1_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_0 = GPA1_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_3 = GPA1_3_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_2 = GPA1_2_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_5 = GPA1_5_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_4 = GPA1_4_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_7 = GPA1_7_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_6 = GPA1_6_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_135 = {_T_128_7,_T_128_6,_T_128_5,_T_128_4,_T_128_3,_T_128_2,_T_128_1,_T_128_0}; // @[CLA.scala 33:46]
  assign _T_128_9 = GPA1_9_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_8 = GPA1_8_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_11 = GPA1_11_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_10 = GPA1_10_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_13 = GPA1_13_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_12 = GPA1_12_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_15 = GPA1_15_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_14 = GPA1_14_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_143 = {_T_128_15,_T_128_14,_T_128_13,_T_128_12,_T_128_11,_T_128_10,_T_128_9,_T_128_8,_T_135}; // @[CLA.scala 33:46]
  assign _T_128_17 = GPA1_17_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_16 = GPA1_16_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_19 = GPA1_19_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_18 = GPA1_18_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_21 = GPA1_21_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_20 = GPA1_20_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_23 = GPA1_23_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_22 = GPA1_22_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_150 = {_T_128_23,_T_128_22,_T_128_21,_T_128_20,_T_128_19,_T_128_18,_T_128_17,_T_128_16}; // @[CLA.scala 33:46]
  assign _T_128_25 = GPA1_25_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_24 = GPA1_24_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_27 = GPA1_27_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_26 = GPA1_26_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_29 = GPA1_29_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_28 = GPA1_28_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_31 = GPA1_31_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_30 = GPA1_30_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_159 = {_T_128_31,_T_128_30,_T_128_29,_T_128_28,_T_128_27,_T_128_26,_T_128_25,_T_128_24,_T_150,_T_143}; // @[CLA.scala 33:46]
  assign _T_128_33 = GPA1_33_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_32 = GPA1_32_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_35 = GPA1_35_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_34 = GPA1_34_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_37 = GPA1_37_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_36 = GPA1_36_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_39 = GPA1_39_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_38 = GPA1_38_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_166 = {_T_128_39,_T_128_38,_T_128_37,_T_128_36,_T_128_35,_T_128_34,_T_128_33,_T_128_32}; // @[CLA.scala 33:46]
  assign _T_128_41 = GPA1_41_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_40 = GPA1_40_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_43 = GPA1_43_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_42 = GPA1_42_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_45 = GPA1_45_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_44 = GPA1_44_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_47 = GPA1_47_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_46 = GPA1_46_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_174 = {_T_128_47,_T_128_46,_T_128_45,_T_128_44,_T_128_43,_T_128_42,_T_128_41,_T_128_40,_T_166}; // @[CLA.scala 33:46]
  assign _T_128_49 = GPA1_49_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_48 = GPA1_48_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_51 = GPA1_51_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_50 = GPA1_50_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_53 = GPA1_53_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_52 = GPA1_52_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_55 = GPA1_55_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_54 = GPA1_54_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_181 = {_T_128_55,_T_128_54,_T_128_53,_T_128_52,_T_128_51,_T_128_50,_T_128_49,_T_128_48}; // @[CLA.scala 33:46]
  assign _T_128_57 = GPA1_57_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_56 = GPA1_56_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_59 = GPA1_59_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_58 = GPA1_58_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_61 = GPA1_61_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_60 = GPA1_60_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_63 = GPA1_63_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_128_62 = GPA1_62_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_190 = {_T_128_63,_T_128_62,_T_128_61,_T_128_60,_T_128_59,_T_128_58,_T_128_57,_T_128_56,_T_181,_T_174}; // @[CLA.scala 33:46]
  assign _T_192_1 = GPA1_1_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_0 = GPA1_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_3 = GPA1_3_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_2 = GPA1_2_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_5 = GPA1_5_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_4 = GPA1_4_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_7 = GPA1_7_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_6 = GPA1_6_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_199 = {_T_192_7,_T_192_6,_T_192_5,_T_192_4,_T_192_3,_T_192_2,_T_192_1,_T_192_0}; // @[CLA.scala 34:46]
  assign _T_192_9 = GPA1_9_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_8 = GPA1_8_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_11 = GPA1_11_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_10 = GPA1_10_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_13 = GPA1_13_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_12 = GPA1_12_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_15 = GPA1_15_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_14 = GPA1_14_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_207 = {_T_192_15,_T_192_14,_T_192_13,_T_192_12,_T_192_11,_T_192_10,_T_192_9,_T_192_8,_T_199}; // @[CLA.scala 34:46]
  assign _T_192_17 = GPA1_17_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_16 = GPA1_16_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_19 = GPA1_19_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_18 = GPA1_18_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_21 = GPA1_21_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_20 = GPA1_20_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_23 = GPA1_23_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_22 = GPA1_22_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_214 = {_T_192_23,_T_192_22,_T_192_21,_T_192_20,_T_192_19,_T_192_18,_T_192_17,_T_192_16}; // @[CLA.scala 34:46]
  assign _T_192_25 = GPA1_25_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_24 = GPA1_24_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_27 = GPA1_27_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_26 = GPA1_26_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_29 = GPA1_29_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_28 = GPA1_28_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_31 = GPA1_31_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_30 = GPA1_30_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_223 = {_T_192_31,_T_192_30,_T_192_29,_T_192_28,_T_192_27,_T_192_26,_T_192_25,_T_192_24,_T_214,_T_207}; // @[CLA.scala 34:46]
  assign _T_192_33 = GPA1_33_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_32 = GPA1_32_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_35 = GPA1_35_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_34 = GPA1_34_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_37 = GPA1_37_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_36 = GPA1_36_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_39 = GPA1_39_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_38 = GPA1_38_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_230 = {_T_192_39,_T_192_38,_T_192_37,_T_192_36,_T_192_35,_T_192_34,_T_192_33,_T_192_32}; // @[CLA.scala 34:46]
  assign _T_192_41 = GPA1_41_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_40 = GPA1_40_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_43 = GPA1_43_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_42 = GPA1_42_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_45 = GPA1_45_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_44 = GPA1_44_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_47 = GPA1_47_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_46 = GPA1_46_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_238 = {_T_192_47,_T_192_46,_T_192_45,_T_192_44,_T_192_43,_T_192_42,_T_192_41,_T_192_40,_T_230}; // @[CLA.scala 34:46]
  assign _T_192_49 = GPA1_49_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_48 = GPA1_48_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_51 = GPA1_51_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_50 = GPA1_50_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_53 = GPA1_53_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_52 = GPA1_52_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_55 = GPA1_55_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_54 = GPA1_54_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_245 = {_T_192_55,_T_192_54,_T_192_53,_T_192_52,_T_192_51,_T_192_50,_T_192_49,_T_192_48}; // @[CLA.scala 34:46]
  assign _T_192_57 = GPA1_57_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_56 = GPA1_56_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_59 = GPA1_59_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_58 = GPA1_58_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_61 = GPA1_61_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_60 = GPA1_60_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_63 = GPA1_63_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_192_62 = GPA1_62_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_254 = {_T_192_63,_T_192_62,_T_192_61,_T_192_60,_T_192_59,_T_192_58,_T_192_57,_T_192_56,_T_245,_T_238}; // @[CLA.scala 34:46]
  assign s_bit_0 = io_cin ^ GPA1_io_p; // @[CLA.scala 41:14]
  assign _T_256 = CLG_io_c[0]; // @[CLA.scala 43:12]
  assign s_bit_1 = _T_256 ^ GPA1_1_io_p; // @[CLA.scala 43:22]
  assign _T_257 = CLG_io_c[1]; // @[CLA.scala 43:12]
  assign s_bit_2 = _T_257 ^ GPA1_2_io_p; // @[CLA.scala 43:22]
  assign _T_258 = CLG_io_c[2]; // @[CLA.scala 43:12]
  assign s_bit_3 = _T_258 ^ GPA1_3_io_p; // @[CLA.scala 43:22]
  assign _T_259 = CLG_io_c[3]; // @[CLA.scala 43:12]
  assign s_bit_4 = _T_259 ^ GPA1_4_io_p; // @[CLA.scala 43:22]
  assign _T_260 = CLG_io_c[4]; // @[CLA.scala 43:12]
  assign s_bit_5 = _T_260 ^ GPA1_5_io_p; // @[CLA.scala 43:22]
  assign _T_261 = CLG_io_c[5]; // @[CLA.scala 43:12]
  assign s_bit_6 = _T_261 ^ GPA1_6_io_p; // @[CLA.scala 43:22]
  assign _T_262 = CLG_io_c[6]; // @[CLA.scala 43:12]
  assign s_bit_7 = _T_262 ^ GPA1_7_io_p; // @[CLA.scala 43:22]
  assign _T_263 = CLG_io_c[7]; // @[CLA.scala 43:12]
  assign s_bit_8 = _T_263 ^ GPA1_8_io_p; // @[CLA.scala 43:22]
  assign _T_264 = CLG_io_c[8]; // @[CLA.scala 43:12]
  assign s_bit_9 = _T_264 ^ GPA1_9_io_p; // @[CLA.scala 43:22]
  assign _T_265 = CLG_io_c[9]; // @[CLA.scala 43:12]
  assign s_bit_10 = _T_265 ^ GPA1_10_io_p; // @[CLA.scala 43:22]
  assign _T_266 = CLG_io_c[10]; // @[CLA.scala 43:12]
  assign s_bit_11 = _T_266 ^ GPA1_11_io_p; // @[CLA.scala 43:22]
  assign _T_267 = CLG_io_c[11]; // @[CLA.scala 43:12]
  assign s_bit_12 = _T_267 ^ GPA1_12_io_p; // @[CLA.scala 43:22]
  assign _T_268 = CLG_io_c[12]; // @[CLA.scala 43:12]
  assign s_bit_13 = _T_268 ^ GPA1_13_io_p; // @[CLA.scala 43:22]
  assign _T_269 = CLG_io_c[13]; // @[CLA.scala 43:12]
  assign s_bit_14 = _T_269 ^ GPA1_14_io_p; // @[CLA.scala 43:22]
  assign _T_270 = CLG_io_c[14]; // @[CLA.scala 43:12]
  assign s_bit_15 = _T_270 ^ GPA1_15_io_p; // @[CLA.scala 43:22]
  assign _T_271 = CLG_io_c[15]; // @[CLA.scala 43:12]
  assign s_bit_16 = _T_271 ^ GPA1_16_io_p; // @[CLA.scala 43:22]
  assign _T_272 = CLG_io_c[16]; // @[CLA.scala 43:12]
  assign s_bit_17 = _T_272 ^ GPA1_17_io_p; // @[CLA.scala 43:22]
  assign _T_273 = CLG_io_c[17]; // @[CLA.scala 43:12]
  assign s_bit_18 = _T_273 ^ GPA1_18_io_p; // @[CLA.scala 43:22]
  assign _T_274 = CLG_io_c[18]; // @[CLA.scala 43:12]
  assign s_bit_19 = _T_274 ^ GPA1_19_io_p; // @[CLA.scala 43:22]
  assign _T_275 = CLG_io_c[19]; // @[CLA.scala 43:12]
  assign s_bit_20 = _T_275 ^ GPA1_20_io_p; // @[CLA.scala 43:22]
  assign _T_276 = CLG_io_c[20]; // @[CLA.scala 43:12]
  assign s_bit_21 = _T_276 ^ GPA1_21_io_p; // @[CLA.scala 43:22]
  assign _T_277 = CLG_io_c[21]; // @[CLA.scala 43:12]
  assign s_bit_22 = _T_277 ^ GPA1_22_io_p; // @[CLA.scala 43:22]
  assign _T_278 = CLG_io_c[22]; // @[CLA.scala 43:12]
  assign s_bit_23 = _T_278 ^ GPA1_23_io_p; // @[CLA.scala 43:22]
  assign _T_279 = CLG_io_c[23]; // @[CLA.scala 43:12]
  assign s_bit_24 = _T_279 ^ GPA1_24_io_p; // @[CLA.scala 43:22]
  assign _T_280 = CLG_io_c[24]; // @[CLA.scala 43:12]
  assign s_bit_25 = _T_280 ^ GPA1_25_io_p; // @[CLA.scala 43:22]
  assign _T_281 = CLG_io_c[25]; // @[CLA.scala 43:12]
  assign s_bit_26 = _T_281 ^ GPA1_26_io_p; // @[CLA.scala 43:22]
  assign _T_282 = CLG_io_c[26]; // @[CLA.scala 43:12]
  assign s_bit_27 = _T_282 ^ GPA1_27_io_p; // @[CLA.scala 43:22]
  assign _T_283 = CLG_io_c[27]; // @[CLA.scala 43:12]
  assign s_bit_28 = _T_283 ^ GPA1_28_io_p; // @[CLA.scala 43:22]
  assign _T_284 = CLG_io_c[28]; // @[CLA.scala 43:12]
  assign s_bit_29 = _T_284 ^ GPA1_29_io_p; // @[CLA.scala 43:22]
  assign _T_285 = CLG_io_c[29]; // @[CLA.scala 43:12]
  assign s_bit_30 = _T_285 ^ GPA1_30_io_p; // @[CLA.scala 43:22]
  assign _T_286 = CLG_io_c[30]; // @[CLA.scala 43:12]
  assign s_bit_31 = _T_286 ^ GPA1_31_io_p; // @[CLA.scala 43:22]
  assign _T_287 = CLG_io_c[31]; // @[CLA.scala 43:12]
  assign s_bit_32 = _T_287 ^ GPA1_32_io_p; // @[CLA.scala 43:22]
  assign _T_288 = CLG_io_c[32]; // @[CLA.scala 43:12]
  assign s_bit_33 = _T_288 ^ GPA1_33_io_p; // @[CLA.scala 43:22]
  assign _T_289 = CLG_io_c[33]; // @[CLA.scala 43:12]
  assign s_bit_34 = _T_289 ^ GPA1_34_io_p; // @[CLA.scala 43:22]
  assign _T_290 = CLG_io_c[34]; // @[CLA.scala 43:12]
  assign s_bit_35 = _T_290 ^ GPA1_35_io_p; // @[CLA.scala 43:22]
  assign _T_291 = CLG_io_c[35]; // @[CLA.scala 43:12]
  assign s_bit_36 = _T_291 ^ GPA1_36_io_p; // @[CLA.scala 43:22]
  assign _T_292 = CLG_io_c[36]; // @[CLA.scala 43:12]
  assign s_bit_37 = _T_292 ^ GPA1_37_io_p; // @[CLA.scala 43:22]
  assign _T_293 = CLG_io_c[37]; // @[CLA.scala 43:12]
  assign s_bit_38 = _T_293 ^ GPA1_38_io_p; // @[CLA.scala 43:22]
  assign _T_294 = CLG_io_c[38]; // @[CLA.scala 43:12]
  assign s_bit_39 = _T_294 ^ GPA1_39_io_p; // @[CLA.scala 43:22]
  assign _T_295 = CLG_io_c[39]; // @[CLA.scala 43:12]
  assign s_bit_40 = _T_295 ^ GPA1_40_io_p; // @[CLA.scala 43:22]
  assign _T_296 = CLG_io_c[40]; // @[CLA.scala 43:12]
  assign s_bit_41 = _T_296 ^ GPA1_41_io_p; // @[CLA.scala 43:22]
  assign _T_297 = CLG_io_c[41]; // @[CLA.scala 43:12]
  assign s_bit_42 = _T_297 ^ GPA1_42_io_p; // @[CLA.scala 43:22]
  assign _T_298 = CLG_io_c[42]; // @[CLA.scala 43:12]
  assign s_bit_43 = _T_298 ^ GPA1_43_io_p; // @[CLA.scala 43:22]
  assign _T_299 = CLG_io_c[43]; // @[CLA.scala 43:12]
  assign s_bit_44 = _T_299 ^ GPA1_44_io_p; // @[CLA.scala 43:22]
  assign _T_300 = CLG_io_c[44]; // @[CLA.scala 43:12]
  assign s_bit_45 = _T_300 ^ GPA1_45_io_p; // @[CLA.scala 43:22]
  assign _T_301 = CLG_io_c[45]; // @[CLA.scala 43:12]
  assign s_bit_46 = _T_301 ^ GPA1_46_io_p; // @[CLA.scala 43:22]
  assign _T_302 = CLG_io_c[46]; // @[CLA.scala 43:12]
  assign s_bit_47 = _T_302 ^ GPA1_47_io_p; // @[CLA.scala 43:22]
  assign _T_303 = CLG_io_c[47]; // @[CLA.scala 43:12]
  assign s_bit_48 = _T_303 ^ GPA1_48_io_p; // @[CLA.scala 43:22]
  assign _T_304 = CLG_io_c[48]; // @[CLA.scala 43:12]
  assign s_bit_49 = _T_304 ^ GPA1_49_io_p; // @[CLA.scala 43:22]
  assign _T_305 = CLG_io_c[49]; // @[CLA.scala 43:12]
  assign s_bit_50 = _T_305 ^ GPA1_50_io_p; // @[CLA.scala 43:22]
  assign _T_306 = CLG_io_c[50]; // @[CLA.scala 43:12]
  assign s_bit_51 = _T_306 ^ GPA1_51_io_p; // @[CLA.scala 43:22]
  assign _T_307 = CLG_io_c[51]; // @[CLA.scala 43:12]
  assign s_bit_52 = _T_307 ^ GPA1_52_io_p; // @[CLA.scala 43:22]
  assign _T_308 = CLG_io_c[52]; // @[CLA.scala 43:12]
  assign s_bit_53 = _T_308 ^ GPA1_53_io_p; // @[CLA.scala 43:22]
  assign _T_309 = CLG_io_c[53]; // @[CLA.scala 43:12]
  assign s_bit_54 = _T_309 ^ GPA1_54_io_p; // @[CLA.scala 43:22]
  assign _T_310 = CLG_io_c[54]; // @[CLA.scala 43:12]
  assign s_bit_55 = _T_310 ^ GPA1_55_io_p; // @[CLA.scala 43:22]
  assign _T_311 = CLG_io_c[55]; // @[CLA.scala 43:12]
  assign s_bit_56 = _T_311 ^ GPA1_56_io_p; // @[CLA.scala 43:22]
  assign _T_312 = CLG_io_c[56]; // @[CLA.scala 43:12]
  assign s_bit_57 = _T_312 ^ GPA1_57_io_p; // @[CLA.scala 43:22]
  assign _T_313 = CLG_io_c[57]; // @[CLA.scala 43:12]
  assign s_bit_58 = _T_313 ^ GPA1_58_io_p; // @[CLA.scala 43:22]
  assign _T_314 = CLG_io_c[58]; // @[CLA.scala 43:12]
  assign s_bit_59 = _T_314 ^ GPA1_59_io_p; // @[CLA.scala 43:22]
  assign _T_315 = CLG_io_c[59]; // @[CLA.scala 43:12]
  assign s_bit_60 = _T_315 ^ GPA1_60_io_p; // @[CLA.scala 43:22]
  assign _T_316 = CLG_io_c[60]; // @[CLA.scala 43:12]
  assign s_bit_61 = _T_316 ^ GPA1_61_io_p; // @[CLA.scala 43:22]
  assign _T_317 = CLG_io_c[61]; // @[CLA.scala 43:12]
  assign s_bit_62 = _T_317 ^ GPA1_62_io_p; // @[CLA.scala 43:22]
  assign _T_318 = CLG_io_c[62]; // @[CLA.scala 43:12]
  assign s_bit_63 = _T_318 ^ GPA1_63_io_p; // @[CLA.scala 43:22]
  assign _T_326 = {s_bit_7,s_bit_6,s_bit_5,s_bit_4,s_bit_3,s_bit_2,s_bit_1,s_bit_0}; // @[CLA.scala 46:32]
  assign _T_334 = {s_bit_15,s_bit_14,s_bit_13,s_bit_12,s_bit_11,s_bit_10,s_bit_9,s_bit_8,_T_326}; // @[CLA.scala 46:32]
  assign _T_341 = {s_bit_23,s_bit_22,s_bit_21,s_bit_20,s_bit_19,s_bit_18,s_bit_17,s_bit_16}; // @[CLA.scala 46:32]
  assign _T_350 = {s_bit_31,s_bit_30,s_bit_29,s_bit_28,s_bit_27,s_bit_26,s_bit_25,s_bit_24,_T_341,_T_334}; // @[CLA.scala 46:32]
  assign _T_357 = {s_bit_39,s_bit_38,s_bit_37,s_bit_36,s_bit_35,s_bit_34,s_bit_33,s_bit_32}; // @[CLA.scala 46:32]
  assign _T_365 = {s_bit_47,s_bit_46,s_bit_45,s_bit_44,s_bit_43,s_bit_42,s_bit_41,s_bit_40,_T_357}; // @[CLA.scala 46:32]
  assign _T_372 = {s_bit_55,s_bit_54,s_bit_53,s_bit_52,s_bit_51,s_bit_50,s_bit_49,s_bit_48}; // @[CLA.scala 46:32]
  assign _T_381 = {s_bit_63,s_bit_62,s_bit_61,s_bit_60,s_bit_59,s_bit_58,s_bit_57,s_bit_56,_T_372,_T_365}; // @[CLA.scala 46:32]
  assign io_s = {_T_381,_T_350}; // @[CLA.scala 46:8]
  assign io_cout = CLG_io_c[63]; // @[CLA.scala 49:11]
  assign io_G = CLG_io_G; // @[CLA.scala 52:8]
  assign io_A = CLG_io_A; // @[CLA.scala 53:8]
  assign GPA1_io_x = io_x[0]; // @[CLA.scala 26:11]
  assign GPA1_io_y = io_y[0]; // @[CLA.scala 27:11]
  assign GPA1_1_io_x = io_x[1]; // @[CLA.scala 26:11]
  assign GPA1_1_io_y = io_y[1]; // @[CLA.scala 27:11]
  assign GPA1_2_io_x = io_x[2]; // @[CLA.scala 26:11]
  assign GPA1_2_io_y = io_y[2]; // @[CLA.scala 27:11]
  assign GPA1_3_io_x = io_x[3]; // @[CLA.scala 26:11]
  assign GPA1_3_io_y = io_y[3]; // @[CLA.scala 27:11]
  assign GPA1_4_io_x = io_x[4]; // @[CLA.scala 26:11]
  assign GPA1_4_io_y = io_y[4]; // @[CLA.scala 27:11]
  assign GPA1_5_io_x = io_x[5]; // @[CLA.scala 26:11]
  assign GPA1_5_io_y = io_y[5]; // @[CLA.scala 27:11]
  assign GPA1_6_io_x = io_x[6]; // @[CLA.scala 26:11]
  assign GPA1_6_io_y = io_y[6]; // @[CLA.scala 27:11]
  assign GPA1_7_io_x = io_x[7]; // @[CLA.scala 26:11]
  assign GPA1_7_io_y = io_y[7]; // @[CLA.scala 27:11]
  assign GPA1_8_io_x = io_x[8]; // @[CLA.scala 26:11]
  assign GPA1_8_io_y = io_y[8]; // @[CLA.scala 27:11]
  assign GPA1_9_io_x = io_x[9]; // @[CLA.scala 26:11]
  assign GPA1_9_io_y = io_y[9]; // @[CLA.scala 27:11]
  assign GPA1_10_io_x = io_x[10]; // @[CLA.scala 26:11]
  assign GPA1_10_io_y = io_y[10]; // @[CLA.scala 27:11]
  assign GPA1_11_io_x = io_x[11]; // @[CLA.scala 26:11]
  assign GPA1_11_io_y = io_y[11]; // @[CLA.scala 27:11]
  assign GPA1_12_io_x = io_x[12]; // @[CLA.scala 26:11]
  assign GPA1_12_io_y = io_y[12]; // @[CLA.scala 27:11]
  assign GPA1_13_io_x = io_x[13]; // @[CLA.scala 26:11]
  assign GPA1_13_io_y = io_y[13]; // @[CLA.scala 27:11]
  assign GPA1_14_io_x = io_x[14]; // @[CLA.scala 26:11]
  assign GPA1_14_io_y = io_y[14]; // @[CLA.scala 27:11]
  assign GPA1_15_io_x = io_x[15]; // @[CLA.scala 26:11]
  assign GPA1_15_io_y = io_y[15]; // @[CLA.scala 27:11]
  assign GPA1_16_io_x = io_x[16]; // @[CLA.scala 26:11]
  assign GPA1_16_io_y = io_y[16]; // @[CLA.scala 27:11]
  assign GPA1_17_io_x = io_x[17]; // @[CLA.scala 26:11]
  assign GPA1_17_io_y = io_y[17]; // @[CLA.scala 27:11]
  assign GPA1_18_io_x = io_x[18]; // @[CLA.scala 26:11]
  assign GPA1_18_io_y = io_y[18]; // @[CLA.scala 27:11]
  assign GPA1_19_io_x = io_x[19]; // @[CLA.scala 26:11]
  assign GPA1_19_io_y = io_y[19]; // @[CLA.scala 27:11]
  assign GPA1_20_io_x = io_x[20]; // @[CLA.scala 26:11]
  assign GPA1_20_io_y = io_y[20]; // @[CLA.scala 27:11]
  assign GPA1_21_io_x = io_x[21]; // @[CLA.scala 26:11]
  assign GPA1_21_io_y = io_y[21]; // @[CLA.scala 27:11]
  assign GPA1_22_io_x = io_x[22]; // @[CLA.scala 26:11]
  assign GPA1_22_io_y = io_y[22]; // @[CLA.scala 27:11]
  assign GPA1_23_io_x = io_x[23]; // @[CLA.scala 26:11]
  assign GPA1_23_io_y = io_y[23]; // @[CLA.scala 27:11]
  assign GPA1_24_io_x = io_x[24]; // @[CLA.scala 26:11]
  assign GPA1_24_io_y = io_y[24]; // @[CLA.scala 27:11]
  assign GPA1_25_io_x = io_x[25]; // @[CLA.scala 26:11]
  assign GPA1_25_io_y = io_y[25]; // @[CLA.scala 27:11]
  assign GPA1_26_io_x = io_x[26]; // @[CLA.scala 26:11]
  assign GPA1_26_io_y = io_y[26]; // @[CLA.scala 27:11]
  assign GPA1_27_io_x = io_x[27]; // @[CLA.scala 26:11]
  assign GPA1_27_io_y = io_y[27]; // @[CLA.scala 27:11]
  assign GPA1_28_io_x = io_x[28]; // @[CLA.scala 26:11]
  assign GPA1_28_io_y = io_y[28]; // @[CLA.scala 27:11]
  assign GPA1_29_io_x = io_x[29]; // @[CLA.scala 26:11]
  assign GPA1_29_io_y = io_y[29]; // @[CLA.scala 27:11]
  assign GPA1_30_io_x = io_x[30]; // @[CLA.scala 26:11]
  assign GPA1_30_io_y = io_y[30]; // @[CLA.scala 27:11]
  assign GPA1_31_io_x = io_x[31]; // @[CLA.scala 26:11]
  assign GPA1_31_io_y = io_y[31]; // @[CLA.scala 27:11]
  assign GPA1_32_io_x = io_x[32]; // @[CLA.scala 26:11]
  assign GPA1_32_io_y = io_y[32]; // @[CLA.scala 27:11]
  assign GPA1_33_io_x = io_x[33]; // @[CLA.scala 26:11]
  assign GPA1_33_io_y = io_y[33]; // @[CLA.scala 27:11]
  assign GPA1_34_io_x = io_x[34]; // @[CLA.scala 26:11]
  assign GPA1_34_io_y = io_y[34]; // @[CLA.scala 27:11]
  assign GPA1_35_io_x = io_x[35]; // @[CLA.scala 26:11]
  assign GPA1_35_io_y = io_y[35]; // @[CLA.scala 27:11]
  assign GPA1_36_io_x = io_x[36]; // @[CLA.scala 26:11]
  assign GPA1_36_io_y = io_y[36]; // @[CLA.scala 27:11]
  assign GPA1_37_io_x = io_x[37]; // @[CLA.scala 26:11]
  assign GPA1_37_io_y = io_y[37]; // @[CLA.scala 27:11]
  assign GPA1_38_io_x = io_x[38]; // @[CLA.scala 26:11]
  assign GPA1_38_io_y = io_y[38]; // @[CLA.scala 27:11]
  assign GPA1_39_io_x = io_x[39]; // @[CLA.scala 26:11]
  assign GPA1_39_io_y = io_y[39]; // @[CLA.scala 27:11]
  assign GPA1_40_io_x = io_x[40]; // @[CLA.scala 26:11]
  assign GPA1_40_io_y = io_y[40]; // @[CLA.scala 27:11]
  assign GPA1_41_io_x = io_x[41]; // @[CLA.scala 26:11]
  assign GPA1_41_io_y = io_y[41]; // @[CLA.scala 27:11]
  assign GPA1_42_io_x = io_x[42]; // @[CLA.scala 26:11]
  assign GPA1_42_io_y = io_y[42]; // @[CLA.scala 27:11]
  assign GPA1_43_io_x = io_x[43]; // @[CLA.scala 26:11]
  assign GPA1_43_io_y = io_y[43]; // @[CLA.scala 27:11]
  assign GPA1_44_io_x = io_x[44]; // @[CLA.scala 26:11]
  assign GPA1_44_io_y = io_y[44]; // @[CLA.scala 27:11]
  assign GPA1_45_io_x = io_x[45]; // @[CLA.scala 26:11]
  assign GPA1_45_io_y = io_y[45]; // @[CLA.scala 27:11]
  assign GPA1_46_io_x = io_x[46]; // @[CLA.scala 26:11]
  assign GPA1_46_io_y = io_y[46]; // @[CLA.scala 27:11]
  assign GPA1_47_io_x = io_x[47]; // @[CLA.scala 26:11]
  assign GPA1_47_io_y = io_y[47]; // @[CLA.scala 27:11]
  assign GPA1_48_io_x = io_x[48]; // @[CLA.scala 26:11]
  assign GPA1_48_io_y = io_y[48]; // @[CLA.scala 27:11]
  assign GPA1_49_io_x = io_x[49]; // @[CLA.scala 26:11]
  assign GPA1_49_io_y = io_y[49]; // @[CLA.scala 27:11]
  assign GPA1_50_io_x = io_x[50]; // @[CLA.scala 26:11]
  assign GPA1_50_io_y = io_y[50]; // @[CLA.scala 27:11]
  assign GPA1_51_io_x = io_x[51]; // @[CLA.scala 26:11]
  assign GPA1_51_io_y = io_y[51]; // @[CLA.scala 27:11]
  assign GPA1_52_io_x = io_x[52]; // @[CLA.scala 26:11]
  assign GPA1_52_io_y = io_y[52]; // @[CLA.scala 27:11]
  assign GPA1_53_io_x = io_x[53]; // @[CLA.scala 26:11]
  assign GPA1_53_io_y = io_y[53]; // @[CLA.scala 27:11]
  assign GPA1_54_io_x = io_x[54]; // @[CLA.scala 26:11]
  assign GPA1_54_io_y = io_y[54]; // @[CLA.scala 27:11]
  assign GPA1_55_io_x = io_x[55]; // @[CLA.scala 26:11]
  assign GPA1_55_io_y = io_y[55]; // @[CLA.scala 27:11]
  assign GPA1_56_io_x = io_x[56]; // @[CLA.scala 26:11]
  assign GPA1_56_io_y = io_y[56]; // @[CLA.scala 27:11]
  assign GPA1_57_io_x = io_x[57]; // @[CLA.scala 26:11]
  assign GPA1_57_io_y = io_y[57]; // @[CLA.scala 27:11]
  assign GPA1_58_io_x = io_x[58]; // @[CLA.scala 26:11]
  assign GPA1_58_io_y = io_y[58]; // @[CLA.scala 27:11]
  assign GPA1_59_io_x = io_x[59]; // @[CLA.scala 26:11]
  assign GPA1_59_io_y = io_y[59]; // @[CLA.scala 27:11]
  assign GPA1_60_io_x = io_x[60]; // @[CLA.scala 26:11]
  assign GPA1_60_io_y = io_y[60]; // @[CLA.scala 27:11]
  assign GPA1_61_io_x = io_x[61]; // @[CLA.scala 26:11]
  assign GPA1_61_io_y = io_y[61]; // @[CLA.scala 27:11]
  assign GPA1_62_io_x = io_x[62]; // @[CLA.scala 26:11]
  assign GPA1_62_io_y = io_y[62]; // @[CLA.scala 27:11]
  assign GPA1_63_io_x = io_x[63]; // @[CLA.scala 26:11]
  assign GPA1_63_io_y = io_y[63]; // @[CLA.scala 27:11]
  assign CLG_io_g = {_T_190,_T_159}; // @[CLA.scala 33:9]
  assign CLG_io_a = {_T_254,_T_223}; // @[CLA.scala 34:9]
  assign CLG_io_cin = io_cin; // @[CLA.scala 35:11]
endmodule
