module GPA1(
  input   io_x,
  input   io_y,
  output  io_g,
  output  io_p,
  output  io_a
);
  wire  g; // @[GPA1.scala 17:16]
  wire  p; // @[GPA1.scala 18:16]
  assign g = io_x & io_y; // @[GPA1.scala 17:16]
  assign p = io_x ^ io_y; // @[GPA1.scala 18:16]
  assign io_g = io_x & io_y; // @[GPA1.scala 20:8]
  assign io_p = io_x ^ io_y; // @[GPA1.scala 21:8]
  assign io_a = g | p; // @[GPA1.scala 22:8]
endmodule
module CLG(
  input  [31:0] io_g,
  input  [31:0] io_a,
  input         io_cin,
  output [31:0] io_c,
  output        io_G,
  output        io_A
);
  wire  _T; // @[CLG.scala 18:18]
  wire  _T_1; // @[CLG.scala 19:18]
  wire  _T_2; // @[CLG.scala 18:18]
  wire  _T_3; // @[CLG.scala 19:18]
  wire  _T_6; // @[CLG.scala 26:21]
  wire  _T_7; // @[CLG.scala 26:11]
  wire  _T_8; // @[CLG.scala 26:31]
  wire  _T_9; // @[CLG.scala 18:18]
  wire  _T_10; // @[CLG.scala 19:18]
  wire  _T_18; // @[CLG.scala 26:21]
  wire  _T_19; // @[CLG.scala 26:11]
  wire  _T_20; // @[CLG.scala 26:31]
  wire  _T_21; // @[CLG.scala 18:18]
  wire  _T_22; // @[CLG.scala 19:18]
  wire  _T_35; // @[CLG.scala 26:21]
  wire  _T_36; // @[CLG.scala 26:11]
  wire  _T_37; // @[CLG.scala 26:31]
  wire  _T_38; // @[CLG.scala 18:18]
  wire  _T_39; // @[CLG.scala 19:18]
  wire  _T_57; // @[CLG.scala 26:21]
  wire  _T_58; // @[CLG.scala 26:11]
  wire  _T_59; // @[CLG.scala 26:31]
  wire  _T_60; // @[CLG.scala 18:18]
  wire  _T_61; // @[CLG.scala 19:18]
  wire  _T_84; // @[CLG.scala 26:21]
  wire  _T_85; // @[CLG.scala 26:11]
  wire  _T_86; // @[CLG.scala 26:31]
  wire  _T_87; // @[CLG.scala 18:18]
  wire  _T_88; // @[CLG.scala 19:18]
  wire  _T_116; // @[CLG.scala 26:21]
  wire  _T_117; // @[CLG.scala 26:11]
  wire  _T_118; // @[CLG.scala 26:31]
  wire  _T_119; // @[CLG.scala 18:18]
  wire  _T_120; // @[CLG.scala 19:18]
  wire  _T_153; // @[CLG.scala 26:21]
  wire  _T_154; // @[CLG.scala 26:11]
  wire  _T_155; // @[CLG.scala 26:31]
  wire  _T_156; // @[CLG.scala 18:18]
  wire  _T_157; // @[CLG.scala 19:18]
  wire  _T_195; // @[CLG.scala 26:21]
  wire  _T_196; // @[CLG.scala 26:11]
  wire  _T_197; // @[CLG.scala 26:31]
  wire  _T_198; // @[CLG.scala 18:18]
  wire  _T_199; // @[CLG.scala 19:18]
  wire  _T_242; // @[CLG.scala 26:21]
  wire  _T_243; // @[CLG.scala 26:11]
  wire  _T_244; // @[CLG.scala 26:31]
  wire  _T_245; // @[CLG.scala 18:18]
  wire  _T_246; // @[CLG.scala 19:18]
  wire  _T_294; // @[CLG.scala 26:21]
  wire  _T_295; // @[CLG.scala 26:11]
  wire  _T_296; // @[CLG.scala 26:31]
  wire  _T_297; // @[CLG.scala 18:18]
  wire  _T_298; // @[CLG.scala 19:18]
  wire  _T_351; // @[CLG.scala 26:21]
  wire  _T_352; // @[CLG.scala 26:11]
  wire  _T_353; // @[CLG.scala 26:31]
  wire  _T_354; // @[CLG.scala 18:18]
  wire  _T_355; // @[CLG.scala 19:18]
  wire  _T_413; // @[CLG.scala 26:21]
  wire  _T_414; // @[CLG.scala 26:11]
  wire  _T_415; // @[CLG.scala 26:31]
  wire  _T_416; // @[CLG.scala 18:18]
  wire  _T_417; // @[CLG.scala 19:18]
  wire  _T_480; // @[CLG.scala 26:21]
  wire  _T_481; // @[CLG.scala 26:11]
  wire  _T_482; // @[CLG.scala 26:31]
  wire  _T_483; // @[CLG.scala 18:18]
  wire  _T_484; // @[CLG.scala 19:18]
  wire  _T_552; // @[CLG.scala 26:21]
  wire  _T_553; // @[CLG.scala 26:11]
  wire  _T_554; // @[CLG.scala 26:31]
  wire  _T_555; // @[CLG.scala 18:18]
  wire  _T_556; // @[CLG.scala 19:18]
  wire  _T_629; // @[CLG.scala 26:21]
  wire  _T_630; // @[CLG.scala 26:11]
  wire  _T_631; // @[CLG.scala 26:31]
  wire  _T_632; // @[CLG.scala 18:18]
  wire  _T_633; // @[CLG.scala 19:18]
  wire  _T_711; // @[CLG.scala 26:21]
  wire  _T_712; // @[CLG.scala 26:11]
  wire  _T_713; // @[CLG.scala 26:31]
  wire  _T_714; // @[CLG.scala 18:18]
  wire  _T_715; // @[CLG.scala 19:18]
  wire  _T_798; // @[CLG.scala 26:21]
  wire  _T_799; // @[CLG.scala 26:11]
  wire  _T_800; // @[CLG.scala 26:31]
  wire  _T_801; // @[CLG.scala 18:18]
  wire  _T_802; // @[CLG.scala 19:18]
  wire  _T_890; // @[CLG.scala 26:21]
  wire  _T_891; // @[CLG.scala 26:11]
  wire  _T_892; // @[CLG.scala 26:31]
  wire  _T_893; // @[CLG.scala 18:18]
  wire  _T_894; // @[CLG.scala 19:18]
  wire  _T_987; // @[CLG.scala 26:21]
  wire  _T_988; // @[CLG.scala 26:11]
  wire  _T_989; // @[CLG.scala 26:31]
  wire  _T_990; // @[CLG.scala 18:18]
  wire  _T_991; // @[CLG.scala 19:18]
  wire  _T_1089; // @[CLG.scala 26:21]
  wire  _T_1090; // @[CLG.scala 26:11]
  wire  _T_1091; // @[CLG.scala 26:31]
  wire  _T_1092; // @[CLG.scala 18:18]
  wire  _T_1093; // @[CLG.scala 19:18]
  wire  _T_1196; // @[CLG.scala 26:21]
  wire  _T_1197; // @[CLG.scala 26:11]
  wire  _T_1198; // @[CLG.scala 26:31]
  wire  _T_1199; // @[CLG.scala 18:18]
  wire  _T_1200; // @[CLG.scala 19:18]
  wire  _T_1308; // @[CLG.scala 26:21]
  wire  _T_1309; // @[CLG.scala 26:11]
  wire  _T_1310; // @[CLG.scala 26:31]
  wire  _T_1311; // @[CLG.scala 18:18]
  wire  _T_1312; // @[CLG.scala 19:18]
  wire  _T_1425; // @[CLG.scala 26:21]
  wire  _T_1426; // @[CLG.scala 26:11]
  wire  _T_1427; // @[CLG.scala 26:31]
  wire  _T_1428; // @[CLG.scala 18:18]
  wire  _T_1429; // @[CLG.scala 19:18]
  wire  _T_1547; // @[CLG.scala 26:21]
  wire  _T_1548; // @[CLG.scala 26:11]
  wire  _T_1549; // @[CLG.scala 26:31]
  wire  _T_1550; // @[CLG.scala 18:18]
  wire  _T_1551; // @[CLG.scala 19:18]
  wire  _T_1674; // @[CLG.scala 26:21]
  wire  _T_1675; // @[CLG.scala 26:11]
  wire  _T_1676; // @[CLG.scala 26:31]
  wire  _T_1677; // @[CLG.scala 18:18]
  wire  _T_1678; // @[CLG.scala 19:18]
  wire  _T_1806; // @[CLG.scala 26:21]
  wire  _T_1807; // @[CLG.scala 26:11]
  wire  _T_1808; // @[CLG.scala 26:31]
  wire  _T_1809; // @[CLG.scala 18:18]
  wire  _T_1810; // @[CLG.scala 19:18]
  wire  _T_1943; // @[CLG.scala 26:21]
  wire  _T_1944; // @[CLG.scala 26:11]
  wire  _T_1945; // @[CLG.scala 26:31]
  wire  _T_1946; // @[CLG.scala 18:18]
  wire  _T_1947; // @[CLG.scala 19:18]
  wire  _T_2085; // @[CLG.scala 26:21]
  wire  _T_2086; // @[CLG.scala 26:11]
  wire  _T_2087; // @[CLG.scala 26:31]
  wire  _T_2088; // @[CLG.scala 18:18]
  wire  _T_2089; // @[CLG.scala 19:18]
  wire  _T_2232; // @[CLG.scala 26:21]
  wire  _T_2233; // @[CLG.scala 26:11]
  wire  _T_2234; // @[CLG.scala 26:31]
  wire  _T_2235; // @[CLG.scala 18:18]
  wire  _T_2236; // @[CLG.scala 19:18]
  wire  _T_2384; // @[CLG.scala 26:21]
  wire  _T_2385; // @[CLG.scala 26:11]
  wire  _T_2386; // @[CLG.scala 26:31]
  wire  _T_2387; // @[CLG.scala 18:18]
  wire  _T_2388; // @[CLG.scala 19:18]
  wire  _T_2541; // @[CLG.scala 26:21]
  wire  _T_2542; // @[CLG.scala 26:11]
  wire  _T_2543; // @[CLG.scala 26:31]
  wire  _T_2544; // @[CLG.scala 41:22]
  wire  c_bit_0; // @[CLG.scala 41:12]
  wire  _T_2545; // @[CLG.scala 41:22]
  wire  c_bit_1; // @[CLG.scala 41:12]
  wire  _T_2546; // @[CLG.scala 41:22]
  wire  c_bit_2; // @[CLG.scala 41:12]
  wire  _T_2547; // @[CLG.scala 41:22]
  wire  c_bit_3; // @[CLG.scala 41:12]
  wire  _T_2548; // @[CLG.scala 41:22]
  wire  c_bit_4; // @[CLG.scala 41:12]
  wire  _T_2549; // @[CLG.scala 41:22]
  wire  c_bit_5; // @[CLG.scala 41:12]
  wire  _T_2550; // @[CLG.scala 41:22]
  wire  c_bit_6; // @[CLG.scala 41:12]
  wire  _T_2551; // @[CLG.scala 41:22]
  wire  c_bit_7; // @[CLG.scala 41:12]
  wire  _T_2552; // @[CLG.scala 41:22]
  wire  c_bit_8; // @[CLG.scala 41:12]
  wire  _T_2553; // @[CLG.scala 41:22]
  wire  c_bit_9; // @[CLG.scala 41:12]
  wire  _T_2554; // @[CLG.scala 41:22]
  wire  c_bit_10; // @[CLG.scala 41:12]
  wire  _T_2555; // @[CLG.scala 41:22]
  wire  c_bit_11; // @[CLG.scala 41:12]
  wire  _T_2556; // @[CLG.scala 41:22]
  wire  c_bit_12; // @[CLG.scala 41:12]
  wire  _T_2557; // @[CLG.scala 41:22]
  wire  c_bit_13; // @[CLG.scala 41:12]
  wire  _T_2558; // @[CLG.scala 41:22]
  wire  c_bit_14; // @[CLG.scala 41:12]
  wire  _T_2559; // @[CLG.scala 41:22]
  wire  c_bit_15; // @[CLG.scala 41:12]
  wire  _T_2560; // @[CLG.scala 41:22]
  wire  c_bit_16; // @[CLG.scala 41:12]
  wire  _T_2561; // @[CLG.scala 41:22]
  wire  c_bit_17; // @[CLG.scala 41:12]
  wire  _T_2562; // @[CLG.scala 41:22]
  wire  c_bit_18; // @[CLG.scala 41:12]
  wire  _T_2563; // @[CLG.scala 41:22]
  wire  c_bit_19; // @[CLG.scala 41:12]
  wire  _T_2564; // @[CLG.scala 41:22]
  wire  c_bit_20; // @[CLG.scala 41:12]
  wire  _T_2565; // @[CLG.scala 41:22]
  wire  c_bit_21; // @[CLG.scala 41:12]
  wire  _T_2566; // @[CLG.scala 41:22]
  wire  c_bit_22; // @[CLG.scala 41:12]
  wire  _T_2567; // @[CLG.scala 41:22]
  wire  c_bit_23; // @[CLG.scala 41:12]
  wire  _T_2568; // @[CLG.scala 41:22]
  wire  c_bit_24; // @[CLG.scala 41:12]
  wire  _T_2569; // @[CLG.scala 41:22]
  wire  c_bit_25; // @[CLG.scala 41:12]
  wire  _T_2570; // @[CLG.scala 41:22]
  wire  c_bit_26; // @[CLG.scala 41:12]
  wire  _T_2571; // @[CLG.scala 41:22]
  wire  c_bit_27; // @[CLG.scala 41:12]
  wire  _T_2572; // @[CLG.scala 41:22]
  wire  c_bit_28; // @[CLG.scala 41:12]
  wire  _T_2573; // @[CLG.scala 41:22]
  wire  c_bit_29; // @[CLG.scala 41:12]
  wire  _T_2574; // @[CLG.scala 41:22]
  wire  c_bit_30; // @[CLG.scala 41:12]
  wire  _T_2575; // @[CLG.scala 41:22]
  wire  c_bit_31; // @[CLG.scala 41:12]
  wire [7:0] _T_2583; // @[CLG.scala 43:32]
  wire [15:0] _T_2591; // @[CLG.scala 43:32]
  wire [7:0] _T_2598; // @[CLG.scala 43:32]
  wire [15:0] _T_2606; // @[CLG.scala 43:32]
  assign _T = io_g[0]; // @[CLG.scala 18:18]
  assign _T_1 = io_a[0]; // @[CLG.scala 19:18]
  assign _T_2 = io_g[1]; // @[CLG.scala 18:18]
  assign _T_3 = io_a[1]; // @[CLG.scala 19:18]
  assign _T_6 = _T & _T_3; // @[CLG.scala 26:21]
  assign _T_7 = _T_2 | _T_6; // @[CLG.scala 26:11]
  assign _T_8 = _T_3 & _T_1; // @[CLG.scala 26:31]
  assign _T_9 = io_g[2]; // @[CLG.scala 18:18]
  assign _T_10 = io_a[2]; // @[CLG.scala 19:18]
  assign _T_18 = _T_7 & _T_10; // @[CLG.scala 26:21]
  assign _T_19 = _T_9 | _T_18; // @[CLG.scala 26:11]
  assign _T_20 = _T_10 & _T_8; // @[CLG.scala 26:31]
  assign _T_21 = io_g[3]; // @[CLG.scala 18:18]
  assign _T_22 = io_a[3]; // @[CLG.scala 19:18]
  assign _T_35 = _T_19 & _T_22; // @[CLG.scala 26:21]
  assign _T_36 = _T_21 | _T_35; // @[CLG.scala 26:11]
  assign _T_37 = _T_22 & _T_20; // @[CLG.scala 26:31]
  assign _T_38 = io_g[4]; // @[CLG.scala 18:18]
  assign _T_39 = io_a[4]; // @[CLG.scala 19:18]
  assign _T_57 = _T_36 & _T_39; // @[CLG.scala 26:21]
  assign _T_58 = _T_38 | _T_57; // @[CLG.scala 26:11]
  assign _T_59 = _T_39 & _T_37; // @[CLG.scala 26:31]
  assign _T_60 = io_g[5]; // @[CLG.scala 18:18]
  assign _T_61 = io_a[5]; // @[CLG.scala 19:18]
  assign _T_84 = _T_58 & _T_61; // @[CLG.scala 26:21]
  assign _T_85 = _T_60 | _T_84; // @[CLG.scala 26:11]
  assign _T_86 = _T_61 & _T_59; // @[CLG.scala 26:31]
  assign _T_87 = io_g[6]; // @[CLG.scala 18:18]
  assign _T_88 = io_a[6]; // @[CLG.scala 19:18]
  assign _T_116 = _T_85 & _T_88; // @[CLG.scala 26:21]
  assign _T_117 = _T_87 | _T_116; // @[CLG.scala 26:11]
  assign _T_118 = _T_88 & _T_86; // @[CLG.scala 26:31]
  assign _T_119 = io_g[7]; // @[CLG.scala 18:18]
  assign _T_120 = io_a[7]; // @[CLG.scala 19:18]
  assign _T_153 = _T_117 & _T_120; // @[CLG.scala 26:21]
  assign _T_154 = _T_119 | _T_153; // @[CLG.scala 26:11]
  assign _T_155 = _T_120 & _T_118; // @[CLG.scala 26:31]
  assign _T_156 = io_g[8]; // @[CLG.scala 18:18]
  assign _T_157 = io_a[8]; // @[CLG.scala 19:18]
  assign _T_195 = _T_154 & _T_157; // @[CLG.scala 26:21]
  assign _T_196 = _T_156 | _T_195; // @[CLG.scala 26:11]
  assign _T_197 = _T_157 & _T_155; // @[CLG.scala 26:31]
  assign _T_198 = io_g[9]; // @[CLG.scala 18:18]
  assign _T_199 = io_a[9]; // @[CLG.scala 19:18]
  assign _T_242 = _T_196 & _T_199; // @[CLG.scala 26:21]
  assign _T_243 = _T_198 | _T_242; // @[CLG.scala 26:11]
  assign _T_244 = _T_199 & _T_197; // @[CLG.scala 26:31]
  assign _T_245 = io_g[10]; // @[CLG.scala 18:18]
  assign _T_246 = io_a[10]; // @[CLG.scala 19:18]
  assign _T_294 = _T_243 & _T_246; // @[CLG.scala 26:21]
  assign _T_295 = _T_245 | _T_294; // @[CLG.scala 26:11]
  assign _T_296 = _T_246 & _T_244; // @[CLG.scala 26:31]
  assign _T_297 = io_g[11]; // @[CLG.scala 18:18]
  assign _T_298 = io_a[11]; // @[CLG.scala 19:18]
  assign _T_351 = _T_295 & _T_298; // @[CLG.scala 26:21]
  assign _T_352 = _T_297 | _T_351; // @[CLG.scala 26:11]
  assign _T_353 = _T_298 & _T_296; // @[CLG.scala 26:31]
  assign _T_354 = io_g[12]; // @[CLG.scala 18:18]
  assign _T_355 = io_a[12]; // @[CLG.scala 19:18]
  assign _T_413 = _T_352 & _T_355; // @[CLG.scala 26:21]
  assign _T_414 = _T_354 | _T_413; // @[CLG.scala 26:11]
  assign _T_415 = _T_355 & _T_353; // @[CLG.scala 26:31]
  assign _T_416 = io_g[13]; // @[CLG.scala 18:18]
  assign _T_417 = io_a[13]; // @[CLG.scala 19:18]
  assign _T_480 = _T_414 & _T_417; // @[CLG.scala 26:21]
  assign _T_481 = _T_416 | _T_480; // @[CLG.scala 26:11]
  assign _T_482 = _T_417 & _T_415; // @[CLG.scala 26:31]
  assign _T_483 = io_g[14]; // @[CLG.scala 18:18]
  assign _T_484 = io_a[14]; // @[CLG.scala 19:18]
  assign _T_552 = _T_481 & _T_484; // @[CLG.scala 26:21]
  assign _T_553 = _T_483 | _T_552; // @[CLG.scala 26:11]
  assign _T_554 = _T_484 & _T_482; // @[CLG.scala 26:31]
  assign _T_555 = io_g[15]; // @[CLG.scala 18:18]
  assign _T_556 = io_a[15]; // @[CLG.scala 19:18]
  assign _T_629 = _T_553 & _T_556; // @[CLG.scala 26:21]
  assign _T_630 = _T_555 | _T_629; // @[CLG.scala 26:11]
  assign _T_631 = _T_556 & _T_554; // @[CLG.scala 26:31]
  assign _T_632 = io_g[16]; // @[CLG.scala 18:18]
  assign _T_633 = io_a[16]; // @[CLG.scala 19:18]
  assign _T_711 = _T_630 & _T_633; // @[CLG.scala 26:21]
  assign _T_712 = _T_632 | _T_711; // @[CLG.scala 26:11]
  assign _T_713 = _T_633 & _T_631; // @[CLG.scala 26:31]
  assign _T_714 = io_g[17]; // @[CLG.scala 18:18]
  assign _T_715 = io_a[17]; // @[CLG.scala 19:18]
  assign _T_798 = _T_712 & _T_715; // @[CLG.scala 26:21]
  assign _T_799 = _T_714 | _T_798; // @[CLG.scala 26:11]
  assign _T_800 = _T_715 & _T_713; // @[CLG.scala 26:31]
  assign _T_801 = io_g[18]; // @[CLG.scala 18:18]
  assign _T_802 = io_a[18]; // @[CLG.scala 19:18]
  assign _T_890 = _T_799 & _T_802; // @[CLG.scala 26:21]
  assign _T_891 = _T_801 | _T_890; // @[CLG.scala 26:11]
  assign _T_892 = _T_802 & _T_800; // @[CLG.scala 26:31]
  assign _T_893 = io_g[19]; // @[CLG.scala 18:18]
  assign _T_894 = io_a[19]; // @[CLG.scala 19:18]
  assign _T_987 = _T_891 & _T_894; // @[CLG.scala 26:21]
  assign _T_988 = _T_893 | _T_987; // @[CLG.scala 26:11]
  assign _T_989 = _T_894 & _T_892; // @[CLG.scala 26:31]
  assign _T_990 = io_g[20]; // @[CLG.scala 18:18]
  assign _T_991 = io_a[20]; // @[CLG.scala 19:18]
  assign _T_1089 = _T_988 & _T_991; // @[CLG.scala 26:21]
  assign _T_1090 = _T_990 | _T_1089; // @[CLG.scala 26:11]
  assign _T_1091 = _T_991 & _T_989; // @[CLG.scala 26:31]
  assign _T_1092 = io_g[21]; // @[CLG.scala 18:18]
  assign _T_1093 = io_a[21]; // @[CLG.scala 19:18]
  assign _T_1196 = _T_1090 & _T_1093; // @[CLG.scala 26:21]
  assign _T_1197 = _T_1092 | _T_1196; // @[CLG.scala 26:11]
  assign _T_1198 = _T_1093 & _T_1091; // @[CLG.scala 26:31]
  assign _T_1199 = io_g[22]; // @[CLG.scala 18:18]
  assign _T_1200 = io_a[22]; // @[CLG.scala 19:18]
  assign _T_1308 = _T_1197 & _T_1200; // @[CLG.scala 26:21]
  assign _T_1309 = _T_1199 | _T_1308; // @[CLG.scala 26:11]
  assign _T_1310 = _T_1200 & _T_1198; // @[CLG.scala 26:31]
  assign _T_1311 = io_g[23]; // @[CLG.scala 18:18]
  assign _T_1312 = io_a[23]; // @[CLG.scala 19:18]
  assign _T_1425 = _T_1309 & _T_1312; // @[CLG.scala 26:21]
  assign _T_1426 = _T_1311 | _T_1425; // @[CLG.scala 26:11]
  assign _T_1427 = _T_1312 & _T_1310; // @[CLG.scala 26:31]
  assign _T_1428 = io_g[24]; // @[CLG.scala 18:18]
  assign _T_1429 = io_a[24]; // @[CLG.scala 19:18]
  assign _T_1547 = _T_1426 & _T_1429; // @[CLG.scala 26:21]
  assign _T_1548 = _T_1428 | _T_1547; // @[CLG.scala 26:11]
  assign _T_1549 = _T_1429 & _T_1427; // @[CLG.scala 26:31]
  assign _T_1550 = io_g[25]; // @[CLG.scala 18:18]
  assign _T_1551 = io_a[25]; // @[CLG.scala 19:18]
  assign _T_1674 = _T_1548 & _T_1551; // @[CLG.scala 26:21]
  assign _T_1675 = _T_1550 | _T_1674; // @[CLG.scala 26:11]
  assign _T_1676 = _T_1551 & _T_1549; // @[CLG.scala 26:31]
  assign _T_1677 = io_g[26]; // @[CLG.scala 18:18]
  assign _T_1678 = io_a[26]; // @[CLG.scala 19:18]
  assign _T_1806 = _T_1675 & _T_1678; // @[CLG.scala 26:21]
  assign _T_1807 = _T_1677 | _T_1806; // @[CLG.scala 26:11]
  assign _T_1808 = _T_1678 & _T_1676; // @[CLG.scala 26:31]
  assign _T_1809 = io_g[27]; // @[CLG.scala 18:18]
  assign _T_1810 = io_a[27]; // @[CLG.scala 19:18]
  assign _T_1943 = _T_1807 & _T_1810; // @[CLG.scala 26:21]
  assign _T_1944 = _T_1809 | _T_1943; // @[CLG.scala 26:11]
  assign _T_1945 = _T_1810 & _T_1808; // @[CLG.scala 26:31]
  assign _T_1946 = io_g[28]; // @[CLG.scala 18:18]
  assign _T_1947 = io_a[28]; // @[CLG.scala 19:18]
  assign _T_2085 = _T_1944 & _T_1947; // @[CLG.scala 26:21]
  assign _T_2086 = _T_1946 | _T_2085; // @[CLG.scala 26:11]
  assign _T_2087 = _T_1947 & _T_1945; // @[CLG.scala 26:31]
  assign _T_2088 = io_g[29]; // @[CLG.scala 18:18]
  assign _T_2089 = io_a[29]; // @[CLG.scala 19:18]
  assign _T_2232 = _T_2086 & _T_2089; // @[CLG.scala 26:21]
  assign _T_2233 = _T_2088 | _T_2232; // @[CLG.scala 26:11]
  assign _T_2234 = _T_2089 & _T_2087; // @[CLG.scala 26:31]
  assign _T_2235 = io_g[30]; // @[CLG.scala 18:18]
  assign _T_2236 = io_a[30]; // @[CLG.scala 19:18]
  assign _T_2384 = _T_2233 & _T_2236; // @[CLG.scala 26:21]
  assign _T_2385 = _T_2235 | _T_2384; // @[CLG.scala 26:11]
  assign _T_2386 = _T_2236 & _T_2234; // @[CLG.scala 26:31]
  assign _T_2387 = io_g[31]; // @[CLG.scala 18:18]
  assign _T_2388 = io_a[31]; // @[CLG.scala 19:18]
  assign _T_2541 = _T_2385 & _T_2388; // @[CLG.scala 26:21]
  assign _T_2542 = _T_2387 | _T_2541; // @[CLG.scala 26:11]
  assign _T_2543 = _T_2388 & _T_2386; // @[CLG.scala 26:31]
  assign _T_2544 = _T_1 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_0 = _T | _T_2544; // @[CLG.scala 41:12]
  assign _T_2545 = _T_8 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_1 = _T_7 | _T_2545; // @[CLG.scala 41:12]
  assign _T_2546 = _T_20 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_2 = _T_19 | _T_2546; // @[CLG.scala 41:12]
  assign _T_2547 = _T_37 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_3 = _T_36 | _T_2547; // @[CLG.scala 41:12]
  assign _T_2548 = _T_59 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_4 = _T_58 | _T_2548; // @[CLG.scala 41:12]
  assign _T_2549 = _T_86 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_5 = _T_85 | _T_2549; // @[CLG.scala 41:12]
  assign _T_2550 = _T_118 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_6 = _T_117 | _T_2550; // @[CLG.scala 41:12]
  assign _T_2551 = _T_155 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_7 = _T_154 | _T_2551; // @[CLG.scala 41:12]
  assign _T_2552 = _T_197 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_8 = _T_196 | _T_2552; // @[CLG.scala 41:12]
  assign _T_2553 = _T_244 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_9 = _T_243 | _T_2553; // @[CLG.scala 41:12]
  assign _T_2554 = _T_296 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_10 = _T_295 | _T_2554; // @[CLG.scala 41:12]
  assign _T_2555 = _T_353 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_11 = _T_352 | _T_2555; // @[CLG.scala 41:12]
  assign _T_2556 = _T_415 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_12 = _T_414 | _T_2556; // @[CLG.scala 41:12]
  assign _T_2557 = _T_482 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_13 = _T_481 | _T_2557; // @[CLG.scala 41:12]
  assign _T_2558 = _T_554 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_14 = _T_553 | _T_2558; // @[CLG.scala 41:12]
  assign _T_2559 = _T_631 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_15 = _T_630 | _T_2559; // @[CLG.scala 41:12]
  assign _T_2560 = _T_713 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_16 = _T_712 | _T_2560; // @[CLG.scala 41:12]
  assign _T_2561 = _T_800 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_17 = _T_799 | _T_2561; // @[CLG.scala 41:12]
  assign _T_2562 = _T_892 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_18 = _T_891 | _T_2562; // @[CLG.scala 41:12]
  assign _T_2563 = _T_989 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_19 = _T_988 | _T_2563; // @[CLG.scala 41:12]
  assign _T_2564 = _T_1091 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_20 = _T_1090 | _T_2564; // @[CLG.scala 41:12]
  assign _T_2565 = _T_1198 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_21 = _T_1197 | _T_2565; // @[CLG.scala 41:12]
  assign _T_2566 = _T_1310 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_22 = _T_1309 | _T_2566; // @[CLG.scala 41:12]
  assign _T_2567 = _T_1427 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_23 = _T_1426 | _T_2567; // @[CLG.scala 41:12]
  assign _T_2568 = _T_1549 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_24 = _T_1548 | _T_2568; // @[CLG.scala 41:12]
  assign _T_2569 = _T_1676 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_25 = _T_1675 | _T_2569; // @[CLG.scala 41:12]
  assign _T_2570 = _T_1808 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_26 = _T_1807 | _T_2570; // @[CLG.scala 41:12]
  assign _T_2571 = _T_1945 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_27 = _T_1944 | _T_2571; // @[CLG.scala 41:12]
  assign _T_2572 = _T_2087 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_28 = _T_2086 | _T_2572; // @[CLG.scala 41:12]
  assign _T_2573 = _T_2234 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_29 = _T_2233 | _T_2573; // @[CLG.scala 41:12]
  assign _T_2574 = _T_2386 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_30 = _T_2385 | _T_2574; // @[CLG.scala 41:12]
  assign _T_2575 = _T_2543 & io_cin; // @[CLG.scala 41:22]
  assign c_bit_31 = _T_2542 | _T_2575; // @[CLG.scala 41:12]
  assign _T_2583 = {c_bit_7,c_bit_6,c_bit_5,c_bit_4,c_bit_3,c_bit_2,c_bit_1,c_bit_0}; // @[CLG.scala 43:32]
  assign _T_2591 = {c_bit_15,c_bit_14,c_bit_13,c_bit_12,c_bit_11,c_bit_10,c_bit_9,c_bit_8,_T_2583}; // @[CLG.scala 43:32]
  assign _T_2598 = {c_bit_23,c_bit_22,c_bit_21,c_bit_20,c_bit_19,c_bit_18,c_bit_17,c_bit_16}; // @[CLG.scala 43:32]
  assign _T_2606 = {c_bit_31,c_bit_30,c_bit_29,c_bit_28,c_bit_27,c_bit_26,c_bit_25,c_bit_24,_T_2598}; // @[CLG.scala 43:32]
  assign io_c = {_T_2606,_T_2591}; // @[CLG.scala 43:8]
  assign io_G = _T_2387 | _T_2541; // @[CLG.scala 46:8]
  assign io_A = _T_2388 & _T_2386; // @[CLG.scala 47:8]
endmodule
module CLA(
  input         clock,
  input         reset,
  input  [31:0] io_x,
  input  [31:0] io_y,
  input         io_cin,
  output [31:0] io_s,
  output        io_cout,
  output        io_G,
  output        io_A
);
  wire  GPA1_io_x; // @[CLA.scala 25:21]
  wire  GPA1_io_y; // @[CLA.scala 25:21]
  wire  GPA1_io_g; // @[CLA.scala 25:21]
  wire  GPA1_io_p; // @[CLA.scala 25:21]
  wire  GPA1_io_a; // @[CLA.scala 25:21]
  wire  GPA1_1_io_x; // @[CLA.scala 25:21]
  wire  GPA1_1_io_y; // @[CLA.scala 25:21]
  wire  GPA1_1_io_g; // @[CLA.scala 25:21]
  wire  GPA1_1_io_p; // @[CLA.scala 25:21]
  wire  GPA1_1_io_a; // @[CLA.scala 25:21]
  wire  GPA1_2_io_x; // @[CLA.scala 25:21]
  wire  GPA1_2_io_y; // @[CLA.scala 25:21]
  wire  GPA1_2_io_g; // @[CLA.scala 25:21]
  wire  GPA1_2_io_p; // @[CLA.scala 25:21]
  wire  GPA1_2_io_a; // @[CLA.scala 25:21]
  wire  GPA1_3_io_x; // @[CLA.scala 25:21]
  wire  GPA1_3_io_y; // @[CLA.scala 25:21]
  wire  GPA1_3_io_g; // @[CLA.scala 25:21]
  wire  GPA1_3_io_p; // @[CLA.scala 25:21]
  wire  GPA1_3_io_a; // @[CLA.scala 25:21]
  wire  GPA1_4_io_x; // @[CLA.scala 25:21]
  wire  GPA1_4_io_y; // @[CLA.scala 25:21]
  wire  GPA1_4_io_g; // @[CLA.scala 25:21]
  wire  GPA1_4_io_p; // @[CLA.scala 25:21]
  wire  GPA1_4_io_a; // @[CLA.scala 25:21]
  wire  GPA1_5_io_x; // @[CLA.scala 25:21]
  wire  GPA1_5_io_y; // @[CLA.scala 25:21]
  wire  GPA1_5_io_g; // @[CLA.scala 25:21]
  wire  GPA1_5_io_p; // @[CLA.scala 25:21]
  wire  GPA1_5_io_a; // @[CLA.scala 25:21]
  wire  GPA1_6_io_x; // @[CLA.scala 25:21]
  wire  GPA1_6_io_y; // @[CLA.scala 25:21]
  wire  GPA1_6_io_g; // @[CLA.scala 25:21]
  wire  GPA1_6_io_p; // @[CLA.scala 25:21]
  wire  GPA1_6_io_a; // @[CLA.scala 25:21]
  wire  GPA1_7_io_x; // @[CLA.scala 25:21]
  wire  GPA1_7_io_y; // @[CLA.scala 25:21]
  wire  GPA1_7_io_g; // @[CLA.scala 25:21]
  wire  GPA1_7_io_p; // @[CLA.scala 25:21]
  wire  GPA1_7_io_a; // @[CLA.scala 25:21]
  wire  GPA1_8_io_x; // @[CLA.scala 25:21]
  wire  GPA1_8_io_y; // @[CLA.scala 25:21]
  wire  GPA1_8_io_g; // @[CLA.scala 25:21]
  wire  GPA1_8_io_p; // @[CLA.scala 25:21]
  wire  GPA1_8_io_a; // @[CLA.scala 25:21]
  wire  GPA1_9_io_x; // @[CLA.scala 25:21]
  wire  GPA1_9_io_y; // @[CLA.scala 25:21]
  wire  GPA1_9_io_g; // @[CLA.scala 25:21]
  wire  GPA1_9_io_p; // @[CLA.scala 25:21]
  wire  GPA1_9_io_a; // @[CLA.scala 25:21]
  wire  GPA1_10_io_x; // @[CLA.scala 25:21]
  wire  GPA1_10_io_y; // @[CLA.scala 25:21]
  wire  GPA1_10_io_g; // @[CLA.scala 25:21]
  wire  GPA1_10_io_p; // @[CLA.scala 25:21]
  wire  GPA1_10_io_a; // @[CLA.scala 25:21]
  wire  GPA1_11_io_x; // @[CLA.scala 25:21]
  wire  GPA1_11_io_y; // @[CLA.scala 25:21]
  wire  GPA1_11_io_g; // @[CLA.scala 25:21]
  wire  GPA1_11_io_p; // @[CLA.scala 25:21]
  wire  GPA1_11_io_a; // @[CLA.scala 25:21]
  wire  GPA1_12_io_x; // @[CLA.scala 25:21]
  wire  GPA1_12_io_y; // @[CLA.scala 25:21]
  wire  GPA1_12_io_g; // @[CLA.scala 25:21]
  wire  GPA1_12_io_p; // @[CLA.scala 25:21]
  wire  GPA1_12_io_a; // @[CLA.scala 25:21]
  wire  GPA1_13_io_x; // @[CLA.scala 25:21]
  wire  GPA1_13_io_y; // @[CLA.scala 25:21]
  wire  GPA1_13_io_g; // @[CLA.scala 25:21]
  wire  GPA1_13_io_p; // @[CLA.scala 25:21]
  wire  GPA1_13_io_a; // @[CLA.scala 25:21]
  wire  GPA1_14_io_x; // @[CLA.scala 25:21]
  wire  GPA1_14_io_y; // @[CLA.scala 25:21]
  wire  GPA1_14_io_g; // @[CLA.scala 25:21]
  wire  GPA1_14_io_p; // @[CLA.scala 25:21]
  wire  GPA1_14_io_a; // @[CLA.scala 25:21]
  wire  GPA1_15_io_x; // @[CLA.scala 25:21]
  wire  GPA1_15_io_y; // @[CLA.scala 25:21]
  wire  GPA1_15_io_g; // @[CLA.scala 25:21]
  wire  GPA1_15_io_p; // @[CLA.scala 25:21]
  wire  GPA1_15_io_a; // @[CLA.scala 25:21]
  wire  GPA1_16_io_x; // @[CLA.scala 25:21]
  wire  GPA1_16_io_y; // @[CLA.scala 25:21]
  wire  GPA1_16_io_g; // @[CLA.scala 25:21]
  wire  GPA1_16_io_p; // @[CLA.scala 25:21]
  wire  GPA1_16_io_a; // @[CLA.scala 25:21]
  wire  GPA1_17_io_x; // @[CLA.scala 25:21]
  wire  GPA1_17_io_y; // @[CLA.scala 25:21]
  wire  GPA1_17_io_g; // @[CLA.scala 25:21]
  wire  GPA1_17_io_p; // @[CLA.scala 25:21]
  wire  GPA1_17_io_a; // @[CLA.scala 25:21]
  wire  GPA1_18_io_x; // @[CLA.scala 25:21]
  wire  GPA1_18_io_y; // @[CLA.scala 25:21]
  wire  GPA1_18_io_g; // @[CLA.scala 25:21]
  wire  GPA1_18_io_p; // @[CLA.scala 25:21]
  wire  GPA1_18_io_a; // @[CLA.scala 25:21]
  wire  GPA1_19_io_x; // @[CLA.scala 25:21]
  wire  GPA1_19_io_y; // @[CLA.scala 25:21]
  wire  GPA1_19_io_g; // @[CLA.scala 25:21]
  wire  GPA1_19_io_p; // @[CLA.scala 25:21]
  wire  GPA1_19_io_a; // @[CLA.scala 25:21]
  wire  GPA1_20_io_x; // @[CLA.scala 25:21]
  wire  GPA1_20_io_y; // @[CLA.scala 25:21]
  wire  GPA1_20_io_g; // @[CLA.scala 25:21]
  wire  GPA1_20_io_p; // @[CLA.scala 25:21]
  wire  GPA1_20_io_a; // @[CLA.scala 25:21]
  wire  GPA1_21_io_x; // @[CLA.scala 25:21]
  wire  GPA1_21_io_y; // @[CLA.scala 25:21]
  wire  GPA1_21_io_g; // @[CLA.scala 25:21]
  wire  GPA1_21_io_p; // @[CLA.scala 25:21]
  wire  GPA1_21_io_a; // @[CLA.scala 25:21]
  wire  GPA1_22_io_x; // @[CLA.scala 25:21]
  wire  GPA1_22_io_y; // @[CLA.scala 25:21]
  wire  GPA1_22_io_g; // @[CLA.scala 25:21]
  wire  GPA1_22_io_p; // @[CLA.scala 25:21]
  wire  GPA1_22_io_a; // @[CLA.scala 25:21]
  wire  GPA1_23_io_x; // @[CLA.scala 25:21]
  wire  GPA1_23_io_y; // @[CLA.scala 25:21]
  wire  GPA1_23_io_g; // @[CLA.scala 25:21]
  wire  GPA1_23_io_p; // @[CLA.scala 25:21]
  wire  GPA1_23_io_a; // @[CLA.scala 25:21]
  wire  GPA1_24_io_x; // @[CLA.scala 25:21]
  wire  GPA1_24_io_y; // @[CLA.scala 25:21]
  wire  GPA1_24_io_g; // @[CLA.scala 25:21]
  wire  GPA1_24_io_p; // @[CLA.scala 25:21]
  wire  GPA1_24_io_a; // @[CLA.scala 25:21]
  wire  GPA1_25_io_x; // @[CLA.scala 25:21]
  wire  GPA1_25_io_y; // @[CLA.scala 25:21]
  wire  GPA1_25_io_g; // @[CLA.scala 25:21]
  wire  GPA1_25_io_p; // @[CLA.scala 25:21]
  wire  GPA1_25_io_a; // @[CLA.scala 25:21]
  wire  GPA1_26_io_x; // @[CLA.scala 25:21]
  wire  GPA1_26_io_y; // @[CLA.scala 25:21]
  wire  GPA1_26_io_g; // @[CLA.scala 25:21]
  wire  GPA1_26_io_p; // @[CLA.scala 25:21]
  wire  GPA1_26_io_a; // @[CLA.scala 25:21]
  wire  GPA1_27_io_x; // @[CLA.scala 25:21]
  wire  GPA1_27_io_y; // @[CLA.scala 25:21]
  wire  GPA1_27_io_g; // @[CLA.scala 25:21]
  wire  GPA1_27_io_p; // @[CLA.scala 25:21]
  wire  GPA1_27_io_a; // @[CLA.scala 25:21]
  wire  GPA1_28_io_x; // @[CLA.scala 25:21]
  wire  GPA1_28_io_y; // @[CLA.scala 25:21]
  wire  GPA1_28_io_g; // @[CLA.scala 25:21]
  wire  GPA1_28_io_p; // @[CLA.scala 25:21]
  wire  GPA1_28_io_a; // @[CLA.scala 25:21]
  wire  GPA1_29_io_x; // @[CLA.scala 25:21]
  wire  GPA1_29_io_y; // @[CLA.scala 25:21]
  wire  GPA1_29_io_g; // @[CLA.scala 25:21]
  wire  GPA1_29_io_p; // @[CLA.scala 25:21]
  wire  GPA1_29_io_a; // @[CLA.scala 25:21]
  wire  GPA1_30_io_x; // @[CLA.scala 25:21]
  wire  GPA1_30_io_y; // @[CLA.scala 25:21]
  wire  GPA1_30_io_g; // @[CLA.scala 25:21]
  wire  GPA1_30_io_p; // @[CLA.scala 25:21]
  wire  GPA1_30_io_a; // @[CLA.scala 25:21]
  wire  GPA1_31_io_x; // @[CLA.scala 25:21]
  wire  GPA1_31_io_y; // @[CLA.scala 25:21]
  wire  GPA1_31_io_g; // @[CLA.scala 25:21]
  wire  GPA1_31_io_p; // @[CLA.scala 25:21]
  wire  GPA1_31_io_a; // @[CLA.scala 25:21]
  wire [31:0] CLG_io_g; // @[CLA.scala 32:19]
  wire [31:0] CLG_io_a; // @[CLA.scala 32:19]
  wire  CLG_io_cin; // @[CLA.scala 32:19]
  wire [31:0] CLG_io_c; // @[CLA.scala 32:19]
  wire  CLG_io_G; // @[CLA.scala 32:19]
  wire  CLG_io_A; // @[CLA.scala 32:19]
  wire  _T_64_1; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_0; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_3; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_2; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_5; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_4; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_7; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_6; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_71; // @[CLA.scala 33:46]
  wire  _T_64_9; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_8; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_11; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_10; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_13; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_12; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_15; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_14; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [15:0] _T_79; // @[CLA.scala 33:46]
  wire  _T_64_17; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_16; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_19; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_18; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_21; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_20; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_23; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_22; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [7:0] _T_86; // @[CLA.scala 33:46]
  wire  _T_64_25; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_24; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_27; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_26; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_29; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_28; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_31; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire  _T_64_30; // @[CLA.scala 33:19 CLA.scala 33:19]
  wire [15:0] _T_94; // @[CLA.scala 33:46]
  wire  _T_96_1; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_0; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_3; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_2; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_5; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_4; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_7; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_6; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_103; // @[CLA.scala 34:46]
  wire  _T_96_9; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_8; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_11; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_10; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_13; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_12; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_15; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_14; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [15:0] _T_111; // @[CLA.scala 34:46]
  wire  _T_96_17; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_16; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_19; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_18; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_21; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_20; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_23; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_22; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [7:0] _T_118; // @[CLA.scala 34:46]
  wire  _T_96_25; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_24; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_27; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_26; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_29; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_28; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_31; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire  _T_96_30; // @[CLA.scala 34:19 CLA.scala 34:19]
  wire [15:0] _T_126; // @[CLA.scala 34:46]
  wire  s_bit_0; // @[CLA.scala 41:14]
  wire  _T_128; // @[CLA.scala 43:12]
  wire  s_bit_1; // @[CLA.scala 43:22]
  wire  _T_129; // @[CLA.scala 43:12]
  wire  s_bit_2; // @[CLA.scala 43:22]
  wire  _T_130; // @[CLA.scala 43:12]
  wire  s_bit_3; // @[CLA.scala 43:22]
  wire  _T_131; // @[CLA.scala 43:12]
  wire  s_bit_4; // @[CLA.scala 43:22]
  wire  _T_132; // @[CLA.scala 43:12]
  wire  s_bit_5; // @[CLA.scala 43:22]
  wire  _T_133; // @[CLA.scala 43:12]
  wire  s_bit_6; // @[CLA.scala 43:22]
  wire  _T_134; // @[CLA.scala 43:12]
  wire  s_bit_7; // @[CLA.scala 43:22]
  wire  _T_135; // @[CLA.scala 43:12]
  wire  s_bit_8; // @[CLA.scala 43:22]
  wire  _T_136; // @[CLA.scala 43:12]
  wire  s_bit_9; // @[CLA.scala 43:22]
  wire  _T_137; // @[CLA.scala 43:12]
  wire  s_bit_10; // @[CLA.scala 43:22]
  wire  _T_138; // @[CLA.scala 43:12]
  wire  s_bit_11; // @[CLA.scala 43:22]
  wire  _T_139; // @[CLA.scala 43:12]
  wire  s_bit_12; // @[CLA.scala 43:22]
  wire  _T_140; // @[CLA.scala 43:12]
  wire  s_bit_13; // @[CLA.scala 43:22]
  wire  _T_141; // @[CLA.scala 43:12]
  wire  s_bit_14; // @[CLA.scala 43:22]
  wire  _T_142; // @[CLA.scala 43:12]
  wire  s_bit_15; // @[CLA.scala 43:22]
  wire  _T_143; // @[CLA.scala 43:12]
  wire  s_bit_16; // @[CLA.scala 43:22]
  wire  _T_144; // @[CLA.scala 43:12]
  wire  s_bit_17; // @[CLA.scala 43:22]
  wire  _T_145; // @[CLA.scala 43:12]
  wire  s_bit_18; // @[CLA.scala 43:22]
  wire  _T_146; // @[CLA.scala 43:12]
  wire  s_bit_19; // @[CLA.scala 43:22]
  wire  _T_147; // @[CLA.scala 43:12]
  wire  s_bit_20; // @[CLA.scala 43:22]
  wire  _T_148; // @[CLA.scala 43:12]
  wire  s_bit_21; // @[CLA.scala 43:22]
  wire  _T_149; // @[CLA.scala 43:12]
  wire  s_bit_22; // @[CLA.scala 43:22]
  wire  _T_150; // @[CLA.scala 43:12]
  wire  s_bit_23; // @[CLA.scala 43:22]
  wire  _T_151; // @[CLA.scala 43:12]
  wire  s_bit_24; // @[CLA.scala 43:22]
  wire  _T_152; // @[CLA.scala 43:12]
  wire  s_bit_25; // @[CLA.scala 43:22]
  wire  _T_153; // @[CLA.scala 43:12]
  wire  s_bit_26; // @[CLA.scala 43:22]
  wire  _T_154; // @[CLA.scala 43:12]
  wire  s_bit_27; // @[CLA.scala 43:22]
  wire  _T_155; // @[CLA.scala 43:12]
  wire  s_bit_28; // @[CLA.scala 43:22]
  wire  _T_156; // @[CLA.scala 43:12]
  wire  s_bit_29; // @[CLA.scala 43:22]
  wire  _T_157; // @[CLA.scala 43:12]
  wire  s_bit_30; // @[CLA.scala 43:22]
  wire  _T_158; // @[CLA.scala 43:12]
  wire  s_bit_31; // @[CLA.scala 43:22]
  wire [7:0] _T_166; // @[CLA.scala 46:32]
  wire [15:0] _T_174; // @[CLA.scala 46:32]
  wire [7:0] _T_181; // @[CLA.scala 46:32]
  wire [15:0] _T_189; // @[CLA.scala 46:32]
  GPA1 GPA1 ( // @[CLA.scala 25:21]
    .io_x(GPA1_io_x),
    .io_y(GPA1_io_y),
    .io_g(GPA1_io_g),
    .io_p(GPA1_io_p),
    .io_a(GPA1_io_a)
  );
  GPA1 GPA1_1 ( // @[CLA.scala 25:21]
    .io_x(GPA1_1_io_x),
    .io_y(GPA1_1_io_y),
    .io_g(GPA1_1_io_g),
    .io_p(GPA1_1_io_p),
    .io_a(GPA1_1_io_a)
  );
  GPA1 GPA1_2 ( // @[CLA.scala 25:21]
    .io_x(GPA1_2_io_x),
    .io_y(GPA1_2_io_y),
    .io_g(GPA1_2_io_g),
    .io_p(GPA1_2_io_p),
    .io_a(GPA1_2_io_a)
  );
  GPA1 GPA1_3 ( // @[CLA.scala 25:21]
    .io_x(GPA1_3_io_x),
    .io_y(GPA1_3_io_y),
    .io_g(GPA1_3_io_g),
    .io_p(GPA1_3_io_p),
    .io_a(GPA1_3_io_a)
  );
  GPA1 GPA1_4 ( // @[CLA.scala 25:21]
    .io_x(GPA1_4_io_x),
    .io_y(GPA1_4_io_y),
    .io_g(GPA1_4_io_g),
    .io_p(GPA1_4_io_p),
    .io_a(GPA1_4_io_a)
  );
  GPA1 GPA1_5 ( // @[CLA.scala 25:21]
    .io_x(GPA1_5_io_x),
    .io_y(GPA1_5_io_y),
    .io_g(GPA1_5_io_g),
    .io_p(GPA1_5_io_p),
    .io_a(GPA1_5_io_a)
  );
  GPA1 GPA1_6 ( // @[CLA.scala 25:21]
    .io_x(GPA1_6_io_x),
    .io_y(GPA1_6_io_y),
    .io_g(GPA1_6_io_g),
    .io_p(GPA1_6_io_p),
    .io_a(GPA1_6_io_a)
  );
  GPA1 GPA1_7 ( // @[CLA.scala 25:21]
    .io_x(GPA1_7_io_x),
    .io_y(GPA1_7_io_y),
    .io_g(GPA1_7_io_g),
    .io_p(GPA1_7_io_p),
    .io_a(GPA1_7_io_a)
  );
  GPA1 GPA1_8 ( // @[CLA.scala 25:21]
    .io_x(GPA1_8_io_x),
    .io_y(GPA1_8_io_y),
    .io_g(GPA1_8_io_g),
    .io_p(GPA1_8_io_p),
    .io_a(GPA1_8_io_a)
  );
  GPA1 GPA1_9 ( // @[CLA.scala 25:21]
    .io_x(GPA1_9_io_x),
    .io_y(GPA1_9_io_y),
    .io_g(GPA1_9_io_g),
    .io_p(GPA1_9_io_p),
    .io_a(GPA1_9_io_a)
  );
  GPA1 GPA1_10 ( // @[CLA.scala 25:21]
    .io_x(GPA1_10_io_x),
    .io_y(GPA1_10_io_y),
    .io_g(GPA1_10_io_g),
    .io_p(GPA1_10_io_p),
    .io_a(GPA1_10_io_a)
  );
  GPA1 GPA1_11 ( // @[CLA.scala 25:21]
    .io_x(GPA1_11_io_x),
    .io_y(GPA1_11_io_y),
    .io_g(GPA1_11_io_g),
    .io_p(GPA1_11_io_p),
    .io_a(GPA1_11_io_a)
  );
  GPA1 GPA1_12 ( // @[CLA.scala 25:21]
    .io_x(GPA1_12_io_x),
    .io_y(GPA1_12_io_y),
    .io_g(GPA1_12_io_g),
    .io_p(GPA1_12_io_p),
    .io_a(GPA1_12_io_a)
  );
  GPA1 GPA1_13 ( // @[CLA.scala 25:21]
    .io_x(GPA1_13_io_x),
    .io_y(GPA1_13_io_y),
    .io_g(GPA1_13_io_g),
    .io_p(GPA1_13_io_p),
    .io_a(GPA1_13_io_a)
  );
  GPA1 GPA1_14 ( // @[CLA.scala 25:21]
    .io_x(GPA1_14_io_x),
    .io_y(GPA1_14_io_y),
    .io_g(GPA1_14_io_g),
    .io_p(GPA1_14_io_p),
    .io_a(GPA1_14_io_a)
  );
  GPA1 GPA1_15 ( // @[CLA.scala 25:21]
    .io_x(GPA1_15_io_x),
    .io_y(GPA1_15_io_y),
    .io_g(GPA1_15_io_g),
    .io_p(GPA1_15_io_p),
    .io_a(GPA1_15_io_a)
  );
  GPA1 GPA1_16 ( // @[CLA.scala 25:21]
    .io_x(GPA1_16_io_x),
    .io_y(GPA1_16_io_y),
    .io_g(GPA1_16_io_g),
    .io_p(GPA1_16_io_p),
    .io_a(GPA1_16_io_a)
  );
  GPA1 GPA1_17 ( // @[CLA.scala 25:21]
    .io_x(GPA1_17_io_x),
    .io_y(GPA1_17_io_y),
    .io_g(GPA1_17_io_g),
    .io_p(GPA1_17_io_p),
    .io_a(GPA1_17_io_a)
  );
  GPA1 GPA1_18 ( // @[CLA.scala 25:21]
    .io_x(GPA1_18_io_x),
    .io_y(GPA1_18_io_y),
    .io_g(GPA1_18_io_g),
    .io_p(GPA1_18_io_p),
    .io_a(GPA1_18_io_a)
  );
  GPA1 GPA1_19 ( // @[CLA.scala 25:21]
    .io_x(GPA1_19_io_x),
    .io_y(GPA1_19_io_y),
    .io_g(GPA1_19_io_g),
    .io_p(GPA1_19_io_p),
    .io_a(GPA1_19_io_a)
  );
  GPA1 GPA1_20 ( // @[CLA.scala 25:21]
    .io_x(GPA1_20_io_x),
    .io_y(GPA1_20_io_y),
    .io_g(GPA1_20_io_g),
    .io_p(GPA1_20_io_p),
    .io_a(GPA1_20_io_a)
  );
  GPA1 GPA1_21 ( // @[CLA.scala 25:21]
    .io_x(GPA1_21_io_x),
    .io_y(GPA1_21_io_y),
    .io_g(GPA1_21_io_g),
    .io_p(GPA1_21_io_p),
    .io_a(GPA1_21_io_a)
  );
  GPA1 GPA1_22 ( // @[CLA.scala 25:21]
    .io_x(GPA1_22_io_x),
    .io_y(GPA1_22_io_y),
    .io_g(GPA1_22_io_g),
    .io_p(GPA1_22_io_p),
    .io_a(GPA1_22_io_a)
  );
  GPA1 GPA1_23 ( // @[CLA.scala 25:21]
    .io_x(GPA1_23_io_x),
    .io_y(GPA1_23_io_y),
    .io_g(GPA1_23_io_g),
    .io_p(GPA1_23_io_p),
    .io_a(GPA1_23_io_a)
  );
  GPA1 GPA1_24 ( // @[CLA.scala 25:21]
    .io_x(GPA1_24_io_x),
    .io_y(GPA1_24_io_y),
    .io_g(GPA1_24_io_g),
    .io_p(GPA1_24_io_p),
    .io_a(GPA1_24_io_a)
  );
  GPA1 GPA1_25 ( // @[CLA.scala 25:21]
    .io_x(GPA1_25_io_x),
    .io_y(GPA1_25_io_y),
    .io_g(GPA1_25_io_g),
    .io_p(GPA1_25_io_p),
    .io_a(GPA1_25_io_a)
  );
  GPA1 GPA1_26 ( // @[CLA.scala 25:21]
    .io_x(GPA1_26_io_x),
    .io_y(GPA1_26_io_y),
    .io_g(GPA1_26_io_g),
    .io_p(GPA1_26_io_p),
    .io_a(GPA1_26_io_a)
  );
  GPA1 GPA1_27 ( // @[CLA.scala 25:21]
    .io_x(GPA1_27_io_x),
    .io_y(GPA1_27_io_y),
    .io_g(GPA1_27_io_g),
    .io_p(GPA1_27_io_p),
    .io_a(GPA1_27_io_a)
  );
  GPA1 GPA1_28 ( // @[CLA.scala 25:21]
    .io_x(GPA1_28_io_x),
    .io_y(GPA1_28_io_y),
    .io_g(GPA1_28_io_g),
    .io_p(GPA1_28_io_p),
    .io_a(GPA1_28_io_a)
  );
  GPA1 GPA1_29 ( // @[CLA.scala 25:21]
    .io_x(GPA1_29_io_x),
    .io_y(GPA1_29_io_y),
    .io_g(GPA1_29_io_g),
    .io_p(GPA1_29_io_p),
    .io_a(GPA1_29_io_a)
  );
  GPA1 GPA1_30 ( // @[CLA.scala 25:21]
    .io_x(GPA1_30_io_x),
    .io_y(GPA1_30_io_y),
    .io_g(GPA1_30_io_g),
    .io_p(GPA1_30_io_p),
    .io_a(GPA1_30_io_a)
  );
  GPA1 GPA1_31 ( // @[CLA.scala 25:21]
    .io_x(GPA1_31_io_x),
    .io_y(GPA1_31_io_y),
    .io_g(GPA1_31_io_g),
    .io_p(GPA1_31_io_p),
    .io_a(GPA1_31_io_a)
  );
  CLG CLG ( // @[CLA.scala 32:19]
    .io_g(CLG_io_g),
    .io_a(CLG_io_a),
    .io_cin(CLG_io_cin),
    .io_c(CLG_io_c),
    .io_G(CLG_io_G),
    .io_A(CLG_io_A)
  );
  assign _T_64_1 = GPA1_1_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_0 = GPA1_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_3 = GPA1_3_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_2 = GPA1_2_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_5 = GPA1_5_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_4 = GPA1_4_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_7 = GPA1_7_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_6 = GPA1_6_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_71 = {_T_64_7,_T_64_6,_T_64_5,_T_64_4,_T_64_3,_T_64_2,_T_64_1,_T_64_0}; // @[CLA.scala 33:46]
  assign _T_64_9 = GPA1_9_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_8 = GPA1_8_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_11 = GPA1_11_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_10 = GPA1_10_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_13 = GPA1_13_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_12 = GPA1_12_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_15 = GPA1_15_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_14 = GPA1_14_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_79 = {_T_64_15,_T_64_14,_T_64_13,_T_64_12,_T_64_11,_T_64_10,_T_64_9,_T_64_8,_T_71}; // @[CLA.scala 33:46]
  assign _T_64_17 = GPA1_17_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_16 = GPA1_16_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_19 = GPA1_19_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_18 = GPA1_18_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_21 = GPA1_21_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_20 = GPA1_20_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_23 = GPA1_23_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_22 = GPA1_22_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_86 = {_T_64_23,_T_64_22,_T_64_21,_T_64_20,_T_64_19,_T_64_18,_T_64_17,_T_64_16}; // @[CLA.scala 33:46]
  assign _T_64_25 = GPA1_25_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_24 = GPA1_24_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_27 = GPA1_27_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_26 = GPA1_26_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_29 = GPA1_29_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_28 = GPA1_28_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_31 = GPA1_31_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_64_30 = GPA1_30_io_g; // @[CLA.scala 33:19 CLA.scala 33:19]
  assign _T_94 = {_T_64_31,_T_64_30,_T_64_29,_T_64_28,_T_64_27,_T_64_26,_T_64_25,_T_64_24,_T_86}; // @[CLA.scala 33:46]
  assign _T_96_1 = GPA1_1_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_0 = GPA1_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_3 = GPA1_3_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_2 = GPA1_2_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_5 = GPA1_5_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_4 = GPA1_4_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_7 = GPA1_7_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_6 = GPA1_6_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_103 = {_T_96_7,_T_96_6,_T_96_5,_T_96_4,_T_96_3,_T_96_2,_T_96_1,_T_96_0}; // @[CLA.scala 34:46]
  assign _T_96_9 = GPA1_9_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_8 = GPA1_8_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_11 = GPA1_11_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_10 = GPA1_10_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_13 = GPA1_13_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_12 = GPA1_12_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_15 = GPA1_15_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_14 = GPA1_14_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_111 = {_T_96_15,_T_96_14,_T_96_13,_T_96_12,_T_96_11,_T_96_10,_T_96_9,_T_96_8,_T_103}; // @[CLA.scala 34:46]
  assign _T_96_17 = GPA1_17_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_16 = GPA1_16_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_19 = GPA1_19_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_18 = GPA1_18_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_21 = GPA1_21_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_20 = GPA1_20_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_23 = GPA1_23_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_22 = GPA1_22_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_118 = {_T_96_23,_T_96_22,_T_96_21,_T_96_20,_T_96_19,_T_96_18,_T_96_17,_T_96_16}; // @[CLA.scala 34:46]
  assign _T_96_25 = GPA1_25_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_24 = GPA1_24_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_27 = GPA1_27_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_26 = GPA1_26_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_29 = GPA1_29_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_28 = GPA1_28_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_31 = GPA1_31_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_96_30 = GPA1_30_io_a; // @[CLA.scala 34:19 CLA.scala 34:19]
  assign _T_126 = {_T_96_31,_T_96_30,_T_96_29,_T_96_28,_T_96_27,_T_96_26,_T_96_25,_T_96_24,_T_118}; // @[CLA.scala 34:46]
  assign s_bit_0 = io_cin ^ GPA1_io_p; // @[CLA.scala 41:14]
  assign _T_128 = CLG_io_c[0]; // @[CLA.scala 43:12]
  assign s_bit_1 = _T_128 ^ GPA1_1_io_p; // @[CLA.scala 43:22]
  assign _T_129 = CLG_io_c[1]; // @[CLA.scala 43:12]
  assign s_bit_2 = _T_129 ^ GPA1_2_io_p; // @[CLA.scala 43:22]
  assign _T_130 = CLG_io_c[2]; // @[CLA.scala 43:12]
  assign s_bit_3 = _T_130 ^ GPA1_3_io_p; // @[CLA.scala 43:22]
  assign _T_131 = CLG_io_c[3]; // @[CLA.scala 43:12]
  assign s_bit_4 = _T_131 ^ GPA1_4_io_p; // @[CLA.scala 43:22]
  assign _T_132 = CLG_io_c[4]; // @[CLA.scala 43:12]
  assign s_bit_5 = _T_132 ^ GPA1_5_io_p; // @[CLA.scala 43:22]
  assign _T_133 = CLG_io_c[5]; // @[CLA.scala 43:12]
  assign s_bit_6 = _T_133 ^ GPA1_6_io_p; // @[CLA.scala 43:22]
  assign _T_134 = CLG_io_c[6]; // @[CLA.scala 43:12]
  assign s_bit_7 = _T_134 ^ GPA1_7_io_p; // @[CLA.scala 43:22]
  assign _T_135 = CLG_io_c[7]; // @[CLA.scala 43:12]
  assign s_bit_8 = _T_135 ^ GPA1_8_io_p; // @[CLA.scala 43:22]
  assign _T_136 = CLG_io_c[8]; // @[CLA.scala 43:12]
  assign s_bit_9 = _T_136 ^ GPA1_9_io_p; // @[CLA.scala 43:22]
  assign _T_137 = CLG_io_c[9]; // @[CLA.scala 43:12]
  assign s_bit_10 = _T_137 ^ GPA1_10_io_p; // @[CLA.scala 43:22]
  assign _T_138 = CLG_io_c[10]; // @[CLA.scala 43:12]
  assign s_bit_11 = _T_138 ^ GPA1_11_io_p; // @[CLA.scala 43:22]
  assign _T_139 = CLG_io_c[11]; // @[CLA.scala 43:12]
  assign s_bit_12 = _T_139 ^ GPA1_12_io_p; // @[CLA.scala 43:22]
  assign _T_140 = CLG_io_c[12]; // @[CLA.scala 43:12]
  assign s_bit_13 = _T_140 ^ GPA1_13_io_p; // @[CLA.scala 43:22]
  assign _T_141 = CLG_io_c[13]; // @[CLA.scala 43:12]
  assign s_bit_14 = _T_141 ^ GPA1_14_io_p; // @[CLA.scala 43:22]
  assign _T_142 = CLG_io_c[14]; // @[CLA.scala 43:12]
  assign s_bit_15 = _T_142 ^ GPA1_15_io_p; // @[CLA.scala 43:22]
  assign _T_143 = CLG_io_c[15]; // @[CLA.scala 43:12]
  assign s_bit_16 = _T_143 ^ GPA1_16_io_p; // @[CLA.scala 43:22]
  assign _T_144 = CLG_io_c[16]; // @[CLA.scala 43:12]
  assign s_bit_17 = _T_144 ^ GPA1_17_io_p; // @[CLA.scala 43:22]
  assign _T_145 = CLG_io_c[17]; // @[CLA.scala 43:12]
  assign s_bit_18 = _T_145 ^ GPA1_18_io_p; // @[CLA.scala 43:22]
  assign _T_146 = CLG_io_c[18]; // @[CLA.scala 43:12]
  assign s_bit_19 = _T_146 ^ GPA1_19_io_p; // @[CLA.scala 43:22]
  assign _T_147 = CLG_io_c[19]; // @[CLA.scala 43:12]
  assign s_bit_20 = _T_147 ^ GPA1_20_io_p; // @[CLA.scala 43:22]
  assign _T_148 = CLG_io_c[20]; // @[CLA.scala 43:12]
  assign s_bit_21 = _T_148 ^ GPA1_21_io_p; // @[CLA.scala 43:22]
  assign _T_149 = CLG_io_c[21]; // @[CLA.scala 43:12]
  assign s_bit_22 = _T_149 ^ GPA1_22_io_p; // @[CLA.scala 43:22]
  assign _T_150 = CLG_io_c[22]; // @[CLA.scala 43:12]
  assign s_bit_23 = _T_150 ^ GPA1_23_io_p; // @[CLA.scala 43:22]
  assign _T_151 = CLG_io_c[23]; // @[CLA.scala 43:12]
  assign s_bit_24 = _T_151 ^ GPA1_24_io_p; // @[CLA.scala 43:22]
  assign _T_152 = CLG_io_c[24]; // @[CLA.scala 43:12]
  assign s_bit_25 = _T_152 ^ GPA1_25_io_p; // @[CLA.scala 43:22]
  assign _T_153 = CLG_io_c[25]; // @[CLA.scala 43:12]
  assign s_bit_26 = _T_153 ^ GPA1_26_io_p; // @[CLA.scala 43:22]
  assign _T_154 = CLG_io_c[26]; // @[CLA.scala 43:12]
  assign s_bit_27 = _T_154 ^ GPA1_27_io_p; // @[CLA.scala 43:22]
  assign _T_155 = CLG_io_c[27]; // @[CLA.scala 43:12]
  assign s_bit_28 = _T_155 ^ GPA1_28_io_p; // @[CLA.scala 43:22]
  assign _T_156 = CLG_io_c[28]; // @[CLA.scala 43:12]
  assign s_bit_29 = _T_156 ^ GPA1_29_io_p; // @[CLA.scala 43:22]
  assign _T_157 = CLG_io_c[29]; // @[CLA.scala 43:12]
  assign s_bit_30 = _T_157 ^ GPA1_30_io_p; // @[CLA.scala 43:22]
  assign _T_158 = CLG_io_c[30]; // @[CLA.scala 43:12]
  assign s_bit_31 = _T_158 ^ GPA1_31_io_p; // @[CLA.scala 43:22]
  assign _T_166 = {s_bit_7,s_bit_6,s_bit_5,s_bit_4,s_bit_3,s_bit_2,s_bit_1,s_bit_0}; // @[CLA.scala 46:32]
  assign _T_174 = {s_bit_15,s_bit_14,s_bit_13,s_bit_12,s_bit_11,s_bit_10,s_bit_9,s_bit_8,_T_166}; // @[CLA.scala 46:32]
  assign _T_181 = {s_bit_23,s_bit_22,s_bit_21,s_bit_20,s_bit_19,s_bit_18,s_bit_17,s_bit_16}; // @[CLA.scala 46:32]
  assign _T_189 = {s_bit_31,s_bit_30,s_bit_29,s_bit_28,s_bit_27,s_bit_26,s_bit_25,s_bit_24,_T_181}; // @[CLA.scala 46:32]
  assign io_s = {_T_189,_T_174}; // @[CLA.scala 46:8]
  assign io_cout = CLG_io_c[31]; // @[CLA.scala 49:11]
  assign io_G = CLG_io_G; // @[CLA.scala 52:8]
  assign io_A = CLG_io_A; // @[CLA.scala 53:8]
  assign GPA1_io_x = io_x[0]; // @[CLA.scala 26:11]
  assign GPA1_io_y = io_y[0]; // @[CLA.scala 27:11]
  assign GPA1_1_io_x = io_x[1]; // @[CLA.scala 26:11]
  assign GPA1_1_io_y = io_y[1]; // @[CLA.scala 27:11]
  assign GPA1_2_io_x = io_x[2]; // @[CLA.scala 26:11]
  assign GPA1_2_io_y = io_y[2]; // @[CLA.scala 27:11]
  assign GPA1_3_io_x = io_x[3]; // @[CLA.scala 26:11]
  assign GPA1_3_io_y = io_y[3]; // @[CLA.scala 27:11]
  assign GPA1_4_io_x = io_x[4]; // @[CLA.scala 26:11]
  assign GPA1_4_io_y = io_y[4]; // @[CLA.scala 27:11]
  assign GPA1_5_io_x = io_x[5]; // @[CLA.scala 26:11]
  assign GPA1_5_io_y = io_y[5]; // @[CLA.scala 27:11]
  assign GPA1_6_io_x = io_x[6]; // @[CLA.scala 26:11]
  assign GPA1_6_io_y = io_y[6]; // @[CLA.scala 27:11]
  assign GPA1_7_io_x = io_x[7]; // @[CLA.scala 26:11]
  assign GPA1_7_io_y = io_y[7]; // @[CLA.scala 27:11]
  assign GPA1_8_io_x = io_x[8]; // @[CLA.scala 26:11]
  assign GPA1_8_io_y = io_y[8]; // @[CLA.scala 27:11]
  assign GPA1_9_io_x = io_x[9]; // @[CLA.scala 26:11]
  assign GPA1_9_io_y = io_y[9]; // @[CLA.scala 27:11]
  assign GPA1_10_io_x = io_x[10]; // @[CLA.scala 26:11]
  assign GPA1_10_io_y = io_y[10]; // @[CLA.scala 27:11]
  assign GPA1_11_io_x = io_x[11]; // @[CLA.scala 26:11]
  assign GPA1_11_io_y = io_y[11]; // @[CLA.scala 27:11]
  assign GPA1_12_io_x = io_x[12]; // @[CLA.scala 26:11]
  assign GPA1_12_io_y = io_y[12]; // @[CLA.scala 27:11]
  assign GPA1_13_io_x = io_x[13]; // @[CLA.scala 26:11]
  assign GPA1_13_io_y = io_y[13]; // @[CLA.scala 27:11]
  assign GPA1_14_io_x = io_x[14]; // @[CLA.scala 26:11]
  assign GPA1_14_io_y = io_y[14]; // @[CLA.scala 27:11]
  assign GPA1_15_io_x = io_x[15]; // @[CLA.scala 26:11]
  assign GPA1_15_io_y = io_y[15]; // @[CLA.scala 27:11]
  assign GPA1_16_io_x = io_x[16]; // @[CLA.scala 26:11]
  assign GPA1_16_io_y = io_y[16]; // @[CLA.scala 27:11]
  assign GPA1_17_io_x = io_x[17]; // @[CLA.scala 26:11]
  assign GPA1_17_io_y = io_y[17]; // @[CLA.scala 27:11]
  assign GPA1_18_io_x = io_x[18]; // @[CLA.scala 26:11]
  assign GPA1_18_io_y = io_y[18]; // @[CLA.scala 27:11]
  assign GPA1_19_io_x = io_x[19]; // @[CLA.scala 26:11]
  assign GPA1_19_io_y = io_y[19]; // @[CLA.scala 27:11]
  assign GPA1_20_io_x = io_x[20]; // @[CLA.scala 26:11]
  assign GPA1_20_io_y = io_y[20]; // @[CLA.scala 27:11]
  assign GPA1_21_io_x = io_x[21]; // @[CLA.scala 26:11]
  assign GPA1_21_io_y = io_y[21]; // @[CLA.scala 27:11]
  assign GPA1_22_io_x = io_x[22]; // @[CLA.scala 26:11]
  assign GPA1_22_io_y = io_y[22]; // @[CLA.scala 27:11]
  assign GPA1_23_io_x = io_x[23]; // @[CLA.scala 26:11]
  assign GPA1_23_io_y = io_y[23]; // @[CLA.scala 27:11]
  assign GPA1_24_io_x = io_x[24]; // @[CLA.scala 26:11]
  assign GPA1_24_io_y = io_y[24]; // @[CLA.scala 27:11]
  assign GPA1_25_io_x = io_x[25]; // @[CLA.scala 26:11]
  assign GPA1_25_io_y = io_y[25]; // @[CLA.scala 27:11]
  assign GPA1_26_io_x = io_x[26]; // @[CLA.scala 26:11]
  assign GPA1_26_io_y = io_y[26]; // @[CLA.scala 27:11]
  assign GPA1_27_io_x = io_x[27]; // @[CLA.scala 26:11]
  assign GPA1_27_io_y = io_y[27]; // @[CLA.scala 27:11]
  assign GPA1_28_io_x = io_x[28]; // @[CLA.scala 26:11]
  assign GPA1_28_io_y = io_y[28]; // @[CLA.scala 27:11]
  assign GPA1_29_io_x = io_x[29]; // @[CLA.scala 26:11]
  assign GPA1_29_io_y = io_y[29]; // @[CLA.scala 27:11]
  assign GPA1_30_io_x = io_x[30]; // @[CLA.scala 26:11]
  assign GPA1_30_io_y = io_y[30]; // @[CLA.scala 27:11]
  assign GPA1_31_io_x = io_x[31]; // @[CLA.scala 26:11]
  assign GPA1_31_io_y = io_y[31]; // @[CLA.scala 27:11]
  assign CLG_io_g = {_T_94,_T_79}; // @[CLA.scala 33:9]
  assign CLG_io_a = {_T_126,_T_111}; // @[CLA.scala 34:9]
  assign CLG_io_cin = io_cin; // @[CLA.scala 35:11]
endmodule
